XlxV64EB    fa00    1f70ܘ)	�b*%�����iڡ��$}�L>�2@�R�o��<$��X%cɉK%k:K��u��D�A�aP�Xu&6��0}�EsV'� "�
kb��BwW�q��X��7&Q�J�����? R���_g��/�`�����b�7ۢ5�3 ���
�Fr �\\8�4���O��Q�9N�%��n��m.�p��<�L��vݚ�f�FT�5�*)�DZQdIՑx#�>v�Uh���A�N�9ߝ�1��_�Y�N�\�fr�U�|���S:xQ`^`	S��:H�g�Q�F��_+b��ҏ4�|ft	!s������mJ0K	��z$�?䇏�G$����yP�%���ݚ {%y8F}�P�B$�܏HȱY���f�):������!)�K�h0�a^���:[m\���a�����E�����*��R<�ꤋ�T�巟@�Lr}Y�	�"���v��^���v|�Hn�M�G������RCz����
h��ȑ��Z_Z�8u4�C�����a�c-A#��^3~�ĽwLuH.��ם ۟�<g�:S/@��<��{�:�{�%lݪEߠ�f,�1��&����4�GA,/�t°�tUtٗ����ʆ��HgB*fi�!��$7ᩧ����PjѶ]��¼�HCܨ�C��Yˢ�z)x�sc��h���� &>�E���E��\�C����J:�%|����}�1><��X�u�����5a�g�sb�ԃé���j�t�P�U�uQ�WjW��-�>��=�����J���h������� ���4��K<#��-R��[h�F�s���xx~�ǡ�$IJ� r�	b{R�dQ4{W���&�[o�aT�B�2�Q��B���SpC`�VDw�F:i�<.C��p؏���$���]�jT�	���zX��&ߝ\v]�W8���4	5GW�2J��=��s�#�
�o$�^�N�h�;~�����5�A���>#7�C-����Z�D8�f���pE\>�"dN9��䯓Q����}��-FK��D��%vxK����x��{~�<a�̞�6��&��{�A�t���A��BY�Y�\���`y��M�Ⱦ�Yv��OUL��$�?x����o��l勖#�H�~�@2b�j,W5�R6$OqxW� ���q����M/Tr��q�#2�b�b���!���m��V��ʦo���P���iiŽ�hO%zs�����[l��9�XY�O"�-����%�弓��j-ɬ�Z�1�'`,����Ɫ� ���;���=0hM|q�
�jt�g�������s�P���WSUX������[��ww����҆��߰��9 nvΩ�d�`5�0B��]�<�f������t8z�&`�����)L	�=���s��� ���Â�s��8�s8%����T.��~k�I��j�a��\�q0�|����:§D��T��PU����4�t+}�KK:��K��e�c�W���Z]�Q�4�Q�~â�L�~����
=^���� ���� %EC+�����p��T"�2���k
Ϡ���$ovI��b��d�j�"���'����������^@�$-���^.V�m�T��@���H�W��2��0����`�|�_v,�B�����_���e�Ω�3y�yHWx~�{uFeg�F��\��gB�}dC{�"���VO3�:[����O�#S�_���"dw��ڨ?5��毶zͶ�H�]"�Q��ce�c�k�'���H�})x����m3M�jܭw)ǈT$B���q�و�j3�JMY1�^��R�(f�V�쫇�8���#@�p}�ng`�Y���g�I�^�a^>�^���4����r��O0}�т9�8���p
CeZ�6�F�33� >��$`�J�X�k���3Ŕ��������cٲ;gGH��V�$�����4���0�wvs�32��{�i�~�j���r�G�;t�M|Jf��!�@�`Ԣ����n%����$#�f~��DgZ�����J�ٸ�6qa��<�i�qD�^3�P�J�� '�	������j)z���u������ڪ�	F�|�
n���G�x��o���1Py��Z������œ���H%FF����&��R �����Ht��Zx���:��2�~��f�C��>��T3���2�6���E-SG��ݍ��&�D{�<�@^q����F�	Xʸ�#&�_,�S7�3!��h��u�P�v�df�ߘ���X����_l��ao��`��B����hpd�� �wxh�G�u�쀞siI4�:�ĵ�\(K�?u��Z���@q(�A���-듙�e��9d�Ra4�Eua�}k��z�@����q��$�|��ږ"��LP�#|��}�A�;�l�M��gf�Q@F����ÚyY��[��/b��m��-�	&2�1(�6>S�)Z���O�T/b-7��i�����Sc����jp����P�[n�� b���ZCDn�0�~�/��U�z0ܧ��ArZwjC2!�#*�o(�jn��
_<��栧��^�7�z����X��7��I@VW.�U(�a��m,7c��q�P-�����&f�-�^$�遷�m��p��鬧��:ɿ$��}�GI�P�ϒ��.�Th%Q��XO\ފ���R�vz#�H��0d:��}ܵ�)�_D k�=$�p��tv�$��k#�"��L�*�O�y�cu	��iV&>�s��Wv��Ea�<�荴ov�"#�=s��;�{��nC�m*�]~� ��,�r�V:|��nA��R�┼����ȿp[���}��vw/�e�Vi=��⬽���fm�m�q4R�����uU�U�`e��K�lC0���#�?��-:;"sX��a�,F�-4̎�o�땊������$�i�A��5��9�~ 
9C��!��N-�-p��60��cQp��m_�L��k�V�<QŽ̦�Y�0��d�-l"b��Eټ�85����m��գ��3C�D�P^���L��eڬ�pf�f-�:�@��`�;+��V����Z2�+���ب��K3Vy#	���$Pq��Q����j�~f��\�_�Ӄ=���0����-�J��]y���K��2�3�j�$"�����M��I�]v`���[�}���X�{�1ά�8�=e=z�˞�m��J������lG}�7)kkH���gO~D%��^�}�����+�P7s{_�D��]-L�Y���;����k���y��&4�F�w&����Kgk�|r�^)�&��$�)�9�4�xVR��Mu�����jA*�׺�X���qL��OE�z�Y�x��͟�KA�������s;�⚪7��� �y�U���'�,͏�"�ޔ݀�Yݱ���<4R�*� �O����M�<�q#��P�p3��2S����+^�X_�4��a����2��=K>�[�*�#�5��P�K���O�˒0anO��bu�xB�s�'�Fp*��,������1��kL�a�XU�Cv�Ҥ��:�5Z*[6]ɜ�~���+�����˫��m;���_�����r���>���9Ѝ趛��!��(�^�q��/Jp�2��cz?�  � V��b�D��ȓ�@#p�RK�&��m��G��j�NIHb�Q�>�~�J"�q�^W�_���� p���B��!�w�-��=Ҹ�������8tZ.��I�mk	��@�̤��1�
� ��&��i� 7^KR6�*��9kZ�����Arn9f�\����hJe��`�D.A�
 ��8s�X�-�=�A�2.y� *+�	��~*�l�Had�Vli�78�_��91JR���G��8�b]PŎ�3/Aޚ�"4s�G��O<�����K�$%+j�wg�8:a� E�T�ΙI�DS���66�������Ebٰ:����簾����!�n�?���2<�|��K.�1��o�-G6E����"̜��^[+��Ҡ�ܖ�N��>agx�Y& �6�������A�Y �A��!�h'u���"�oq�$%��?���I�T](���h���3��o;(t�G��:I�=\UԮ��E>n0���X�:7�����l�⑳a��pVZF�]�-X���4��{9��;���	��):�j��)��w{���j���)��(�̭C��p���5c	���Ҋ��lr�lժ�1��� �í�(�b΄��r���!F�<Y"�{4;��=�J�w��˽̜���-W����Ń���nh=n,��r�L�miθ�y?l�4p����>���*7g4Eq�D��sk���th��?biec����U͸Y��_��tu�4X�%>�s�B����`#P���j�]˚�W�կ1�a��[�ۭ�^'�p��2h�6��M���s��;�D
�NB66��&�8,�����vl���!'S�̂#���	!EƼo����d+�]�b�-�zE�,��6t�_-ԨV��6�����`&�����}�eb�YՎ��s�Jl�mx3��ͳ��A2����fg<G�k��
��)�t�pߋ'����yv| �˚��^>Z�1/V��Ƅ���^-�/B��Vý�_m/����QCFk��`�l#���ߖ�E)���a�Ѥ����R)e����#����Ά��Ш8;��4 U�"# S���ٟ�͑;�7���XQ�����	�(q�,2T+��r*����4<�U�v�/��J{y�f��{聇�e�t���09�>ż��nH�s�i�!k�3(�j����܋g�{��!9���|�r�)6i��_Y(gk��R���x#S!����w�߂Q����O��y�J��zC��Ѳ�-菬><	����&뎣׶�w�{�9(�[��i�q��zlu�����$s�V�}X��h,~t�xx��͠���E�A��TSɼ���N���H�vz�f)�z*F ����G;t��[��/M������g��'sg�gr��M?hU\%9�ܭ�i�Ҷ�D��ap��2_m��X�F}��uW0�������1��?��%�7L�b���R�D�a�K �Lne�W��Huv	����bȕ��r<B%�]�Ol��B�R1g����)�G��pmp]��wDڭ�[M�k�E�1%�JB��4��F2��|v�j"�љ����2�^d;�;���d-2�u5��? O(��[��pù�'�7�����S/����=(�e��T�8x? ��e�=�;��:BakzeCy�w�ǟ���v͘�{��	�A�b�R��gI��Q�S�y�L-x�i"x��Ğ���U�Μr��m� ��~1�r0!��s��ޗ��)��d3t3-�ќ=�zECEt��u����qF����[�M:h�NQ�tnt���FxƵ�p�fQ'��g��#�BǶ'Q���@_�/ztS����XԢR�ᗁ��:m�\s��޸���UY=^��qβj�z(��G�+*��U����#�܆]V�i�L�L-+�����8�L'�F��23#�y�\݋�|�螺eud�ӾUC�/�}������;UЕ�>Zqv�V2y����TŤ$���U2�5���snw%�e�ۨ�/,-���ğ�\�ޣ|}�@�����	�����7�O��.���z���Z�h�>�~mSD���J~z��T�4b"��7�>W��E��9��b<�z�y���+'��q9�=I�z�[�F�Y��B��+{j�����Z Ű����3vX�+�/r�DL�-iQ��<Hd7:N���۶j0嚨8hJ;�hI��=���2pq |��B�����J�q�N�o�`sсRIo0O|z��%k�K������gu)�t2�3����L����å5 t��s�Z�Kx`k
��ɳ���j��轐�u����vif ��br�K�=����@���I4R�JY}S�.ÿ,�kȿݧYj.�"tA����|+�,~*����K�g|k�c)��p��J��K~����Y�w.�d9y��j`��J`<�
�Ix�v�����f�c�.�B�*�ࢩ�}IH��1c0�3ٱ�L\C�\<��ے)Y�oy8�Ո��L$X2'�N�a`a�\Ŏf̑֞R]a �J5�;KM�_�ե���mm�"�������jRiu����ȌKΤ�eW���B�z0%;74��Z��н�8���\��l�~�DJ=e���c�2!A�|�O0�0}�":SAGN�7|[��f�T%8-�5BŇJ�8��*�)`#�;��B,�~��Rˮ�r��ʓ͖��I�}��EGx��f�fj1P�j����h��]a(bz�7c��[���ݔ����?<H��x�����ר?g�E����0�7���(I֟��?E�Cn��{>z:�� �P�l23�G�yo�����,RT+�s���gG�����.��cy��g�K��TdԑH�߅�r�M���U3�1Hv�L�����0�=p��n/�6��w��o��ͦ��t$s)�K�IF��g�U��6i�@C�IC��� ��a��\�(���2,|�Ȁ�T�8��v��r�j��s]!�8��!��&�w���0���7��n�	̹�I�IͶ�ǅW-����I�VL���<��i��+a4��8��T��~�=���O�B3+WY����݋ɤ4.�Z��|6D��e���pY�w���0
�*��Re�1���E�y�v�D��|z �qv\���Vx���)��׸���׋:�%�����C���&���Q�y�����i ��#�"(��r	���-C����硫 ��3$N�=�ǟ�7��B�I]?�,���;�ڟ�M��ᰃ�J����� �&%�<�e0׋m�P?��H0Dr@%�x�L̘v�r��7K��S�ډG�n&x%����揽�|}�u�}|���1\# .��L��p8XѶW�	}����7�b����$tuס����3��3����k��`��Ȁ+8�jW�U��g��b�zoZM�Pck��Var��;��[��QE���+mg ����ae�
P�>w`��Fxu:�"����df�Է8�|`� .h0�"sb�CQ������T6�@��E�㑾�K%���j�~/���8y6���v{��Jt�Kzl���7�rJYD2>A��?�砧����]�40ߌ?��w���I�V�ٟ��Mq����M~�� >�Ƿ���@)��mL��� �_�1�>/�41�Q�j)R��9Q�����ђ� ��y��Y��&�8s��^{�~)���NP�;�Fe���|�_����o�Uf̭���.�����'���ƛN��M�h:��3���N�y��C�ܚ�?�:3��n"g�q�	��H��dnH�H��C.�/z��@)�i�|Y ;݅���)�6�g�3�\^CKt�c�M�|O�Sܹ��u���TO<���K�10Dۯ�N{m҆h���(��	����f��(���2fS�E&b���|GH�G<�g�>�*�CM7��=��)���Ӓ�9k�kG�^����ݖz' �G2����!�F������l�����T�VugC�f]9�,�蛏[��r:3�C𘹗��}�=�۽�QI0��v����"��U�n�,(`X�����,n�s���d�'!�CޭtQ�.�5ͬH]��b���{��-��]CXLx����oG�I������p�o��&���L��`�AR���I�]����H d�۞K�y����>�
P�ķS=���Rb�v'aZ~��.��t�$˰�BU�y��يT��ÀY)VY��	�e;�-r��-��+���ܗYd��&�E]Ծ��n�
+g��JOz��6���8<�%>8)�9a�ƍ!hsEֆ�Ы�T�Ѕ����1�+�#-�$2b!.6�n/���#?��u,�8%rH�7���
�
���ujw=7Rft5dP�XlxV64EB    fa00    10c0O��}:�3��f�(��
���#�Y��1Xy��;P]�9>��V�0T�[^^�Y����E�$�^�٭��-��2`�y��n���ι��H�y�詵ϖt��˼��V%]b9�2�3��r���,�$E0�����¸�t��:e���!!�h<^<��d �ڇ�r9c"W�;��|�����6�l��j;4|o$ձ�� z����\r��\����t�g{���`�?؛��Y
�>ݕ/����tN��I���CA�������B.H� @�smJh��n���e-��@�X��I��ϋ��É����i��qr4����\�H+�a��h����_�a��p�[k��/X�����Blgq!wJ�f�h�i_�p��aK4������ 2�����\����Z7g[(�4��|D5X�ge5��H�B�\*��(���ǟ�^g1 k5�Bd�m�j�T�x®p|*��-����f���n����Sx��[��'�0UחX�� �&�o۱�u�Qq睿o�딐A���hkºƊםL0ҍ�)'5��ΰ��p��J�@i`aE���BW��Z���K����}õ4�4����� G=�ed-T߂F�6����!��C����u6�GB�_<I)��GȐ���</�b9f��LF/��L�����F7�hC
D�@+TC����	<� �V��Ӏ��e�8$�����f�43a>�@�L�.3함�W�[~Pb�dc�-a�4�4�zOT��Y?ܖ9x>h���1�E7�L�Ԛ�m�eG:1��F���^_4�s�#j��v�_?��\�Ӳfy��Y�#�ݟ]e�hn1�B�/�n�6ܜ�f����}4��8�ܬ�LFg@���g�����|�,����?��$���tx`��5�'����0�q����k�!E��0�RͼL��߹>iS�i��5��J��u>Ww'!�-�����QŚ�� � p�[���!��
bw�k�5����k��FZ�lnŀXc���^v���
�(RPnJ颿�4�-��v� ��>7}ޤ������q|���/��TpJ�i��o�fx�F	�d{��G%m-�R��E/k����Z��A<�RE�+S��Zk�����җ�y�=,3\�,�o͏Z�ꖉ���^T�vG�Tϥ�{�%h顖H������Z\�����,Qlo�a'H{������v�N�o=����_���pJ¢�:F�"�U�s+�" ��
����F_�"�9��>�#�q��u%�Qg"�Փ�E�'��_�����i�b>٪��␬9��6�;�������t��UD���ZH��b�j9^���S ���r�I�3i.�@�����b�����1���_u������C��O({���j��fw��7:�n�n�!WFY���wz~/�0݆-�5�>RK�2�����ٖ��I�W��X�mSIO7�{�'G�s�4|�����^�g9�A��"�G��Y�@j�Ʋ���۰�ϴ�sK�k������*��l[2:�	��q���0�7?���['�Ε`���^����O�@������	�)oȹ�=,1nˋ�$��%"L�d�He��b�_�a��Lv@�/�� +�o]D�G����^�h$��ΠǓ`�g�9�^K[�!訑�$�DWb��D
�4ւH�"0K �PnXu�V��k���ε�/���rw���� y�5�J5�eNb�)�gG�N�M����L>P�F�������T��� T�<e���?�;�#V���)��TꗞC4�&����tO�G%�?Y7�Eǁ�g�;ʊs�K~�;)~�@&{���S W�H�pc����W�κ��ʹJ�Вݺ��5I�~�HxI�.�"5�M�VSN�SQ|F����c~y,�{OA�
�#�o\>k,�+�B�2�xC��ry�Z�(R��rA�R�X-l����N"�9�Z]Ч���p�<�0_�Wqn3�Лҫ��c��냶�rҷ�˷�Ą˜���d2dP9dp���1��Fͳ��>�A^��� 4Q��f�r��[Y��z&U���� �Q9�	�!)E�8�K�e�l��2en
���i	�N�T��$��&��A%�!-y�\W!ꯨ-t����7D��$��-MZ�ib�°�K��SO<���eq���w�i�5Pw�!ax`q8��
����lo<i@�D���u�JĻ��ƴ8�y!%�3�*�tҗ���6�O�_Z<� ����dm�ߋۤd�DM�W�z&���ͤi���|�rk��-��Fj�׮Μ�-���Z��d��0k_6�y{�ְ�9���1���ǀ���%��mF�2��w����{�4���P����%�vc� Q>|,|�m��d{.��7и�)q�W�%�W��m�CD f�9 [o����]͛{G�7�?���gM����y�$�C�x�K�Ǆm�/t���?�w�"����\��`��ڒ��6My$��6�4+���u'I-��	TƂ��ʉ��{Ǝ����mE+q��k[���2���ٞ�)+Ǩ���dWA�2��Lz!�01��q;%3A��:�uDK�u�+:�����҈��v/֌#E��v�m���tm&<m�u"^�?	J�%>.��M#ȭu��h�]`r��y����0�-�S���Q�j�ʷ�P�3�[��@�W��#c�uF~��FP�H!~���dAw��	�퇳��-A��+2�c
���sN>92�Za��5|t,����T��(��$��!S�3|N����Wڞp�_`�7�I*>�4\ �n�OjR,��I�L��RE�臋��	�b[�X7z�|����"�Z��B�P ���A�$2�q$�ě�@����g���AN�:a�R5�I+�V�X�0��0����#�;z��u�Rµ5������0����|���	�z8LH���^+>ƿ�'.�� �3q�.rH�N8�	<�2<�9��+~��� ����w'9���K��/f�%�x/M��s��m�E�q�MբP�#�C�X�
�ʏ����vb��9���ڽ�5be@�w��Y�n��'8�}n��,�L������������j}��5��7�8ԙum+p;�lA|��3���ҝ��qi�{��LpP$۽%V6;._�~S��\X�>M�5K�\�h,^���"��8&�>q�E��Ӎ�/��Y穃0��Z�JѹR�}�/;V�	I��P4�RH?�'���f~K!�cݕf|�g�+8&�:�OJ���L�2m��nLX�>򙵍�w�����x��m��-�*�d�����̨�aU����0�䑏�gE;ϕ�3�m���־K��{%��# 1�<2���4l�A������3��sz&+`��IY�[�<y��h��Ԅ$�Ī����8�#"l�DY,}i�U�:�rM�+���4Ձ�4)U:f��үpӑ�1�.�ٶBِe��
A���1'P��a������$�4b�'���@x43�ޑ\�7��w����'��ȣ�qj��m�ÄI�����½;ˮ�*l鲠��h7��zV���.���Bs�	����^�]G�V��[��&_�O�kccr�g(�zZ�4��E ����a��̒~�"� �{�J��wC�ƪ�(8�q �)��`wR���365�k#�����V\:�����я�{�	7q-�B~�@3��$�3qh�� �Ը�ɫڌ<�m��N��P�#� �����ݘ��"��yDf	�����u,�Z�˦ss� 1�+M�޻���`��M�I��Zg2U+�����$庑zPy6��j�u�y�!]$kQJ���*hm��[�T��z&�v!;��qY���'�+��G����R:�Xov�=�ư�k&:��&�茪���zgg&)������	�� �7�U�gc@� ������ݩ\݈%�ZA��h�2^̜��؊:������(Z���LIRk�Q���k�nX�Q�:�g�T��d% �����n%mIm�i�u5g��v�,NE�f\�&f���{_<DR�M�E�/X�?b�i+/��dT�z_�\A_�f�p��CF8�&�����<jɧ�6�XO)B���Z��R3�&(��mo��U�w�}�/zn���$���J)S�`:��m�|p\>��n���,
,��γ �����|�Z��=�G��1y���@��)������"�@�ml�e��|�΄q����OSҊH��ţ��XlxV64EB    fa00    1140[.�PjX����;�M�D�������x�\��i��46���bUqS	򮣲�?�/�A�`��1�S� ��)�<u�.jd�cG<���v \w>ۜK�W��,������@��\�4�/j�+�ɴGI�X���T�.P�Ӱ�L�q��,��""&9�P��n���1!��!�8&L:˟߮7c��u��=�Ih/���/0�����U�i�K�W\�N�'�{�ڥ_o���V�R��B��� � ���6�MQC�E��䌺�5��g��:�+�m�ݓ4"��劓R�b�K���(�߀/`omq�/bɤ+�k��s�P"+�Nя����G 2�M�7�M,���4�y@.aTX��;�X"<Eҍ0\��Xt>$L��ڸ���QI����W��譧��1�2�B'��\�k4L������p���������z��W��+vά��o�����MYp9�t?�ܧ!̟  �"N�M	<i0���m������0��$X�;�V?�+�aѦ�LxJ~�g6-����R<�ah��60�Уۖ�EH\)�HM�R7�"�x��-mir�Qd8x����f@񦜂�@���Ǫ��9P=��K�7�ӓT�>�׋�-�W�W0R�S
0��;1�MR���u#���ঘt��o����L��x��H+6��?���> .�?Lg��3�$�)�P�p���I�n9x�����6_��ѣ�(�4P��)��Q��`^=W;&��^�ԋ"']��a��qE��kk��m����묹���木���[���W���myL���h:��VC	�@l��U(n��m�%B�JZ/S��#��9�x�8X����#����`���6��������:4�����@�m�,�	gj���W6�'�K����P4��?4� ���n?�!oP�R��)H��u���^$@]k�i�!�h�!�Y�ȇ�m�ŭ5$d�� 6%�g�N���O�PE.���r�T�2�}��p��A:$[|�L��N��L�A�DX.�z�s�5AI�jR�)�L-o=n�ˮ"�4��OwbVYL�2�1y$�(r�ц��İ/����q�T�`��5��f�����N�⎹+� �����:B��5Q���/�Fw\$�2#�67P�;(�"Z�n=�,��2�f��e����ي�*d8cʃ�|���7�l�2��L���&����;��r�va�o�Q&H��y�8|,�Q+1)�����j�l��S���p�IGb&���
���yahN�aS��K^�|=
k�H�J�(��A�񄅋�g��w�ʰN���Y�(��Ɓ�3�T0��ZP���:���~�T�K-�ZN��R���ۦIE�G����ѱ���^6�~�g{	ӈ����F��j�?�s<?�*0����h�P{,Vo����ԜJ�ڲ�gi�h�=����f������I��J��dc��d������(��Q�64�[[�V�_H;Wp�]�X={-Kg3TYf͜J�w������'�!�R�Y��3�D��∓��i9�&���KqN��@w`G���
|{�Ёgu(s�'��6�0maJ�%��5C�iA��}��w�=pN��pT�6;�i��ΌO�H�v��n���?P9=���/�4U�� <�U_�M��'��cp���A�i����4�p]ܖ�ȭI������a�2��Y��������B?�@��}�L����������9���OP�T�5��&��T�p�A�[�/ غV\��'D{��W�=3�y�NB�*n%��#$!y��]T����<���F�-!i	է�z	���=y[OL}X�r��tf���?(/r#{x��E7�Y(*>��/�i4(r�U*E�ֆr�M^�}%�]�8D2:Ԓ��>�F3|�8w��R�bM��6�#�rW&�+�������$$5	�0�����
X���8]9f�����������:ގ��=�!�I�1���о���q��Pf�cc����O�t�&k&nw�aeb8y�dWj�wC=���Bo�����n��M�M�X��{�u�E�QlS��\I[�x}�ze!���≸��?�������V�p�|��������$���w�}lj�M��B@3H�X�F}�b���`��d#�W�3� �Fc@����U�v�U�fK���G�����cD�O�=�����6�'�B�y����)Fz����G�)7�:N��F�L��I����`�'���#'ۗ4Ĝ����`�O�B~�M�O�t�ҧCa�y�{+	A�2�j�'��\ q�ք�&���@�D��x'BN�)j̘��{�Қ!:�t�#}�($h*�1��o�LEMaa��H"���`�@?j<'g��׈�Y��c�*s#�81�veBnʪ]�y�{��ݪk�v*�M��h��}���RW�P���������p��c�/E�G�M�:�Tc�$�Q�JO��w��M�)��=��o\|�E�>w=\%���"Bf<�x�ǽ��a��5�tQ�Go���H��M%�.,�)�7����p��rn�X8����g�x:7����«M���㲸}D5����Gv�la����8k��jT-��U�g��A5j��%8unP�K{Y]sC/BƘ߶�؄i�d���|���+(��`㚬Z=�S5Y��،8TB��E`�K]�G�q���O���{*�;]�� y֛�v��c��gM�
��w��Ɖ���񊒮���|�p
�BamF���k��N$8̽7	ݙ*7���<m lc�xWc<Ʊ7�"a�sVoTS�ib��B�:�/��8J��$��>�:3*l8����;?��P��q&�$�Ⱥ���+ن�5���f��]�PJ��
���v:�2�^�$7Jy�vqi�ưA��(?�yl�\��f@:w[.TL�z`v���"�=k�j7C���ǁ�r��I �����xy�]Dw�i��('��>Sn0 �J�F�+#d<��N�{t���t]n���QZK���\8�v�9�����%P�@%�(�y+���I
#�`Y�hG��"C���[�20(�8T��ۺ�P�`
�D�^g�P��htI�����	m�d<���O�W�q�@��>�1�R���Ѝ�;��ԣ�����W�ë7H!�e ��� B�_y��-��v7�la^\jp�D`B%��Y=��	v��ن֛�ǧ�l�CU��V��u�z/#q&� ��I������iq��|.���쐭�� ������������"Ǩ��ܚ\�)o�%��$���{���(�Eb�n�3
z`�����"�����4TG�鱁��U��ǧ5��a���@��T�fT"j���j �6�@�^0q&&�v�(6m�Q�!�	�a�s�ݴ$f�������w+�>'Ϣҥ��qK��r_j+���5�,`�ҍ�k�좒������C�뎿��G����t��:��^�歓��A�~<�l]3�z��hH��b�9$�� �DѰ��A���d��'�6�ʔ�gUTF�3�]����O@K�¹�{=~o�3�-��e5L��Մ���'�.���>�)�| >m�HwIp��c�јB6Yp9ǫk��N�˱k%+��=�RF���<�޷Vy۳Զ3^sY1�z�w�t1����ؔ��%��N�J^	B��>� %K�?��3щ��ds�([,W�?KE�}��
��Њ� 諒0^�z�Y%��0��'��Yot���m*�*& ���Bçz�ؕs䯭ۅ)��_ ����(pcux�Q�E]�����~X6��`zY����`�d��nf�	�B>��=}�5^��8y�){�XRA�g8(� ]�1�}
�A�FK�������E���4Of�,H���nƂ�^��}���=���c�X�9PD�p��@��ai�0Z�Vu�k=�e!�;߸E�8�l�˂N�$y��U ��O~�2+�ٕG�� �?aG�O�p�:��x�䃙�P��9ׁv�̅�ȱK��MnX�b��󓘯���ea���"��`��4	Q(���ɀ���jr �/���x��u��=Ո:�I�$y�/i�:�	]�@wz�#������շ����&���%�î�FiȌ�˶	�r��@@��0���ղT����{N�$�ѭ�|/�C�����t��Q�Y#f0��� �4�S�+��4�g4���jz�N9��F��
L�.S������d�'|��aX���}��'�`*������I�U��|ʬ���:��D�=�:����H�Iȗ�=���-I9g�e:�W��ł��V�z���.C)�MMpe��t�1�c�����)~�x?�\3��SG����v^���p&�
V���y�XlxV64EB    fa00    12e0�^����m��,��EVy�ͩ*���ٽ�<�u��8shH�h����[3�+��� 	�x'�
C�����>���nB)_�Pa�|�i��)<.~���i��t�i��H�('Kl^=
��Q�f�
C�5��q�̄�"���V�@a�=-������䊕����m��5�d�w�s��Jtr(��@�����~y-4%�G�p��\i�����3�΢�,����բ�<~>�D(6�M��Ҽ�ǀ�wO�'�����!�w�G�r��~�O��I&�I�H|��r��~�rҝ1���4A�]�����:s��`x�6�&�!3v3�*a>�'�Vx8'�i�L�J�]�	��J=!��@џ������z��ra�,�0Pݸ�\�P�6��	j'2�fxlvQ"�
K���"- 3A�p���l�Ո:��'�r=�s���iMݧ�>ˑ����o�u΂�?����H�7s��/�;�>�ԛ�s;	}h�� <e �q��9�6���\�����LM�|�i/[#<c9�赲9�պ�fڰx*Х���4�Ϻ*���JJq87��	��f�F����ʥQ��y.�
�}�/���g�ܘ�_#Z5�A���O���p*�c�]�?S�oV�Z>�����D���7��^��$�w�w��/`ߍy��Id��P�%��d���v�0�/��\"ۀU�ɏIm�Ek&T�w_,9�Ϛ�*�,��r��D7��n_� �����lL�\� ԗ��Y3� �q�Q�Z�.�����������M���,��Ž;S<�96} >�=���b��	�L�v�%bow2���
�(�"_��|�~-B;�6CQT�N1;�웻���]�M�����)yLp$� �QY��	���N�$��|�:F�� f�ن�
I����
�LP&=CAV6��3�`�8	��`1���T���1�+�[E���-��{D��^�6H���}��ԸY�sT����^���g����$����W|ń��A�4>����ޖ�$b�z�_�C��K��@��t�T��z��u�����^/����Y@��r�,mD�c��Df�UXFI\x?����k�DFz�.��{��� Ȗ2�>3.��[Mf��(hc�	��{gNn,槯��b7��:v�=<�R��h#���`��v��)�ǎ�*|�d`xo����թ���z�V*ȣGl��N���������A�hZ�H8��a�9�E����d&Q����/�q�(�C����рR�m�"$(5��lP(��~8�q��Hf�}r�H27��� �64��v1�]�0���z��
ou]-��.FwTǄ�x똯���#�S�IѺ�l�%#[@d5Jɸ�@�Î�e)�]锽P����T0ɿ�-�ޤ�&$���L}i���/���.�O�Jgk5}����!�>��˝2>a����9�J�S1#�*� �&L$����˅�o���F�z�u�J�l��I��P5���޵2�}S&�j(][_4	DX����3��� ?�ɂo[����B��RĲ��c+�nײ��Y�3QI�m�V�]-�.����:C.�(  ?���d��2k&b9FeSt&�'ڻ�����S$��͢���$�Ľ�!
�w����|�������'vq�B�5}����|�!�Y��\�ث�A����]��[��'�g���f����9'S�f�n:5�1��j�9�/L����Y[.�k�i
���)Cw\_�p��+ֳ����
�w�4���t��S���j����dLa`��+y��	�{)m6C��M�g�Ra|�T-&]Yä�"�b/Qp�_CUPW�0��/� �O���I�?C\�\򿔤N��[ftp��`Öl��\�19(�5�o'�@}k������oȰ���e��6��)��x�ēa�V�
.���[�Mmڼ�?Z���|){��D: ����9�l��L����h��r����(맛-?�Bbp�����m=)?8�BV��T��Ar��~���l�?���;�_�f ���֖���{�f�C�?,���zd�?�ޭ�Ci�"C�c*�h�EO~���{d>(�zj�ٗ�½�q��h��*�r#�=���*	�"�#�M����z�������\��;��w�w�E��	��L�N(�8�ɗ<���;4��hq��ddYr�C�iwr���(�TՄJ���t`�tg��1i%�R͹x�1���'�K=�m�� D�\sq����`��d�M��=7­�kmR��x%D8��@[�N��gh�3�R  O��ʭ:Qp���k��u_�H"%+�Y������u�2l��G�0o�*9�o���%<�r�ۘ-#XkbZO��.^��$��S� �c�[��=[
�$a�Nc���'��WsP:sǌ�7%9ZC�OpQ��2{OD#��tw̄5Y˟�\���`u�9+0d�_u�^���%]�����Y,W��&�,��ѱ�g�.��0��"��>��Y"l9"����>P)����>�.^�;���)x��5<���y�'u?q����:�v�t���K��#���p-Fe��>9�G�ۀ�bYM(�.���J}�,�[��$�:�(6`�{�lz�*@vr���h������~�ƫ��h��Ϯ��e���Ц��%WT,��Wz���2�| [|������%��C�(�iK3-vt}��dpa�l�����=w�št(��{MYҚ�
y��ֺ �n[�������D�Ly@�G����ɛ��[ϼل���� �����������7E!PΟQ���hq>(�^��\�Jɮ\�>�����R'p��C���9T�Р�؝y�2>?\�
9��N�`N�g��5Ƭv���0O�sC0 (E�b�c���''��F���(jo���0���X'���|�\'�~�'���ճo��?�b��j�q:�[�/�PRE�b�� -)�<W�;�1�d�����/-o��f��A��Π��@4��]ߟW�cht��.8s����!�^h�����͔]Gz�ǩ�v��	�}S�Y2W�B�0��T�p�6�z�*�f�0�|*糀���/ߩC����=��@Fsůf�)��R��/��<zqȰ6=7$�����_�g��&��9n��-A�u�`���%v	M�(ٖ�k��-��D��b3R( �Q�1��M��L�J����j�Z�#�Wr �i�i�=�ko���MC� [���2���C��v¼��!���Y�����G��.>v���N��E$��F�Z��v0Bp�Y����ind�	�D4��*�]�X�;1�I)S�-t+����f��H��t&�{7\#��t�QUDENiޖN�1�K%?c����,1�\��
�O��8o���|w��4������k��f��XH��S����`��H�Z��$�pU+%���A��m	�?����3�IO��-K꩸�S�\�nѪ�WkNG��t6tNv�cM_X܃��Ne�A�_���L�JlL�<m�D��N����w@��������ʹL����E�����\ �d�W�.�o�)���Ř~�S�5x(���;������r�c/�E��*~7��N5�3-�Ĵ�U�uQ�v:�n�/T
#r*����zi#�A�A0�=�����'p9�:�ۮ�3yVmtN�������,�
����_1d,�O��Y)��mRH>�Ԟ>ذ&�]�4���VnB�5bDg�ǝ�C�ugd}]���v�
��H��:=��{V�dr���ON�)�]m�o``P�徇P��9��#P>�H��K�h_�y�1��0�߽^:U<2m����sG'�3E�̕����NM�j�p� �E��:Q��E_xļ�x(�]�!8p�$�LxD��<22A���[qp�����k��������U]v@��N{�2�_���
��q�x[�%#l��,5�d$�l��w�: *Ļ�e��\�{`M�����	�L�����F���`-!�-�;c��w��Kom��nB]�d�H悔����7�UH<���.{8��GU�u��Q��+���5^2[����"rl�K��6����%dg ֞�[-!Z5xvo�0e�'�he\��Ssj�em�.:Zj���K�"������}�NѤ}���ۥQ4_�陫�6�S?U����-D'"3u��`��i�p1�NtQ��ci����9��#�ĵ>�p��sU	����"dcMhX��ђ}�V[�Dr$�*�j�����#;���~�G�mQ]z���]ӯ��bd|����E����>=_z�%g�(���H���zd�ژU�p�@��r�ÆG��	�Mc��zټ�+i��E��פ	8�j�Z�i8�#�2�+4���1��;���R[-��+�J"f�z��q�ትeBIt{�^:7���-����˦:# 2���Yu�q[B�A`���-0�]������ט�7d�&w�'Y^��7���=oTސzd���^�d4�*S�,�|i⥧��A�6�<�p�$������f'k����8�����#�a\���=�V��(������OËͭP�@���f�!D=��uM{5+k�fA��q�9{J���}Q�Ͻ
VU�{V4��&*с�$�	��
C��έ�6��R4��������6;W���WȐ*lv���B*��E��}��T	�k�I\�T�N�i7����z|7����\ߗ�gM�dDd�A�%�D^p}���<[�{���ZfMw��Ka.DiI1XlxV64EB    fa00     f50����,x�ӝv�E����Z(����Gd�%Hǻ�Јَ��r�\*M�6f8���탘�v(S+��vK�����[��;�
���_ ��B�լC�٢��F8�����^&;Q�-Ot��N=6>�E����%[}�}}�n���fe�o��4���59ǖ��4�~`��	^�H�V��M��|8�Q�����Oyp�n�@�>Sg��	]C`#���9�H������Ի�S������,����9���!%������A�S
O�p��2�T]f��m���`.�VnL���+������)&�r��/����#P4����1����F��z�o��b�8Џ����k��F�T`�л_͕ڪm<�2^�)�C"�7���=)=T닚�/��c	.]Z��z�p�Y�H��ß{'�*�<o�+�E�̎u�-e_��r�ǤX�·�h���Qxn.L,o�]�4U
���S��DN�ow�]���%'X���G��|vQ�W���O~D����Dv`��s%�����K^��!4HG�q5��
�s��w�̒ن�8�(R�ēܹ�ƃ�o~�>�S8��}C�rH�3�o::�~ Y�P���F���W�l�'�������� �w�����]�Z ]�0�z�+�XDq�ȓ��l)X҈p��"U+��l�1I���u!31���6�~$��ހ�a�A��lD����OU�I�S��������y�������&�oO�/V��hd���Q�!���ӊ'q��<D��Q��H$��fB_z�%�I����z��j¼.�v=���i������Lw���0���z�o40�Q���Љ*��M�*��S=@֎�������L�\ͦ�_	�H�R�o��=�t��p��&�Ʋq��S�j�(�K��%/I8�z�0o�&~K�G<�7���H��N�y��a1X�b�ּk3�*HC��[w���o3��5ڏ�9)	3�������?FP�n��9O;I?^�lI�,���� ^7ԥ�!-�������p�x$N�i�$���pM��u�[\��NDEU�8=d�'�d��qʿ�T+h�Ō[���S�?Z�����ٙ��q����/��"��h���C�/��1��+ii���)�>�j�hD/�^e������\_-�����[�@�lB�v�H7��~�?���5�C��a�j����y�@����ԍ��������ov�~H���ݟq?E(;!��P���obu�����Sk����D� m��@|}��O|�|���b�2�>�7��b'�:
/�٧�	�]>%�2KU�OC/�l���WJ�?�K�W�0,��0�F_(�HL�J���U�E�9��,t�oд��a�-��Ag>��l2���K8���6����0`^��j���B��)��6v�RY��F��ʹ�y��Hx���+��y����Ɵ�zB-�(!Tf2KT��|��%[��OfL������Nb���uKN��3�SD`d]x$~�p�̵�ߥ���?�=N<ڮ$��Z�
��J������g@�mYjj%w!�J�/��ڳNIG��a�r-ͤ/�`����v���|�1`p1�hд�����%�k� �����^Fӟ?�����l�N<	��v0��	�C��M}"��-���AUv���8�s���Tz� ���Z��ƚ샥�؟��`a>"P��hȩA�������&kH��"Q�3��ˊ}�Y��헠w�<�I����I ��% �خn睸7�
ŷ1Z�8���#u��}�+,���I�P�U�?���,x2˕>�$�g}LX����v��0H��Y�����!��ٚ��ڡ�2�p0n�� ����#�j�v��T������W�|{b(K���C����I�<�C_ܳ��B��U�ǃ���K��/��Z؀����I۔��+��0�G����A��B��S�˼��,u�R9�}XA����wHGNU�ᮌI �d��4ܟ�����%w�!=�� qN8��j�/S�y�fd9~�8�5�$T��Š� �DoM+��k=IgOmAS�����v�>]�wQ���R�QV��m[���^=G�ưܙ{W.[���]rT2~CK�Xeu�~d�E)Q?9={���N��d��<>0~�����`}��t��R;��m���]�9[�z_��6�Pz	��nR<7��� jZ����=DB�R� �R��x@as٢�>���(�b��������-t�R��^�J��r29��~�@�*K%A��sH�0~Y��A�EY WF�ҭ�ױ���DsB3�:���������n��w�q_˸����;��.���\�V,`]�a��5<\�o��̺��/��݇M�^r�k�6C��~�w����P%׮y���֘kSЖ��^v����/���C�
��J��΢���~�����FR4�8��c���9��͙0������p�T����#k/��å~C�����T�o�IA�t��L�[O\w2^3����F7c0'^��)�T"qq��D]1��NA:!J����'+�Jx\��$E*q�X�h��*��l�02��y��q�ã�sa@�K.�=X�[��hlzY}r�^"�3E�_�%�"F0\BG� �}���� �ZT `UR��T����%��� 0/�϶��u��K��њ���>��d���)�@�*�%a�K6����KHq%r�B��g^(�[�2ǥe���vu[���0�t����dح��	E��]�҂�d�Ԫ>�eM"��7_(<O=3L&�=�t[���*�=Z/8%��/4�'�f���O��AzWVjM�X����������F*Q�Q4��G��[rA��m:紤M8%�s�*�넹�f����Z;�fX���n�����n,�E^rc��m�a�ӹ�9�˫E��L���A�U�ӞM���t����*O�/�7C�Q�s���v������A+��3c�0όI"���}�<H�5���ץZO����^�"*�"����T�8��@�@#�:z����k�U���"H���<n�d�&�ͤ�+B���%�����6&�K��┦�4	��M���N6e��a�a|c��,�'�u����u�x`�v'�����h���59��ln��q���;rl�Dθ�����ѫP��Y�^I�B>�`k�6w>��N,��x��T��a�S����5���� p'fz_���� }QF�m~�9��i�.KJ�fJ~���OLK'[yn�p�
.�h,�%��o`����&k��u �i}���iX`<wm�O��z�,����. '���T}�xYц���,I�vp�� _#��n/��_$���6�Wޏ��*����WY��@`���9 ������8c��|A}M�W��kZ=�E��7^��w���}�h�j�y���6"#ѳ������z���Yk��7���#��3�N	�dq$z���?�V̰~�HY�ixne;]�-�d���H5)�q�`6�Cܼ��'=\7o���2�T s�r���v�YCUH��wyv�v�,���l9VL�(e!V#��-�)�X�m��_3s���
x~u\$V ��s��#
2�bŮ�|"����Z�<.9�����u��QF++���J���Y�ֳ�9���tO�J�-�.�j[��\,��"P�Yn(8�Ꝗ�,�K(pm?G*Ҧz0ƕ%�R}PE�w>A3�<��t�3���菡J���	�7�W깱��~���pБ ����~��C�����叙e0��\�n�^_jX2�� ���P���3Jf�Y�<�kƹ�S��-,lg��
�mEk�lW���^l#�Id�d� ��@�qXlxV64EB    7795     6c0TAr�^S	��E���Q�U�N�* �璌sZE$X�l\lI?����>�)� Y�sT�!T��@XuږE��"Kp�HM��B�M�:A���4�.�I�&��?N����
�Χ{��S\���b��+"7k�&H��f2
�ʝC�D�W�>���6���+j�}x�K��~f��1h;���u�@VU^Lp���c&�n.�4����H�����*͑:<	H�gŅj,=�~��W:����ڨv��Ωͽ;���>�*�^�� �"�k+G� �' 0�?��(�2�?rx�g[���Sm��&TR���V�ڼ.d!f%ѴY��C�lS�b���{��l�����?���~?�̕���N��ugu8B���g{�6 J��<�2Y��i�������b:z�j�3��1F�#���E�fg�*�VF��R�&����9�6�}��^B��WM��d�'���l�;]��7���� �~���G��������RőQ6~W��RE��.�Ϸ~>�r���
cu���q����6����5��-}$=j���`�U��!Sͳk�,E-4�7��jP"@����0��r��Wqr{��nHb	�"�m,�'�[�rzAv���|0v|�����V���C��3S0�+�����"�_��jz�uB�-����i�M��4��$G�%)."�YI��:�MȞ,\����e>��b֤D%�k��iC+��EP�6^���n=��� ���)[*��Gd�b=�Z��[�f��ù�����bil�268j�B�$"t�'3�w��K�����m�~�蚚h�����������c���X
�p�j�2H�/�)�2%|�I��M�L�_�T��O��C�E~L�`/�g=$���!|.롈�����?ԫi*��%>��ס4�*�����W�zG+��f�w"/j�F�+��_VǼ�B)aN���.�8��񞍧1YӧۘLfc6���j�Sl(�4o�ދ��(��q!�U�u��|5��·p#���	_~���\�zs��Ɩ�����&���Ǘ����Ih�X��%տ'I��#�>�?D�����"|���&`њ�$L[U,`��r��ӥ:�vV���f�'R?�ᒕ�(,=Ϫ؟��N���K #�/���Y�|�e���Hi6�jI�Q��u"MwģTfH�9�>�RW��V&��x�)�?�*��+%�ɘ*�yӇ�lR��gݻ	�Ť!��(A�0	F�)!(�{L�gj!(N�	�UD��h�;Y��]���pMR�������&^��pII�͛� ����tEc�{a�h�g�m����%ך��I��(��I��n��33�� ����N���]�#OZ���(�޸$c�Y5������
�7pZ��	d��O&{Yg��$z,h�(���R�+ﵩ�7���\���
�j-�.��$3���l ���A/��J��Lѫ�����K�A>��u=C��Ɇ��.{��ؓTphh`#A���|���Zʨ�cu��j�3�1��֯� �J���,�R��|�Ũ����谖��e�!�O�e��.|�E3P1Bհ�az�U�o3"*��g]��c}�J����vYB ��#�΃KP�����q+�@��?��ک�}T���z�<<j,rU����m��F�`T���2�
�yJ��Cԧ�ɼ�x�oji�