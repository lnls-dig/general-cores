XlxV64EB    2608     9d0\8�e��~��~`KL<_�s�ńӂ#�x�њ�}���?���&��Ú�P��?9�����O��ߛ�����oy�i�~j�t�5f�{�T[���J�Ɓ��$���UA�:�.�(Ji�1u���+����®QŽ�~"��:g �o�ӗ&`�{{�k�2!DO�{��Hy��m�߹��A�~��lMDl@<�#{Z��^��>7)ljr۟��p�~7JT>�獽�	����/���'h���m?C����Q喸���Ὓ^��i��Q��DY��K��ҪoѸ�7�q+&k.���̜i����q�':��n�t�e5l�jsZ�HJL��!\��囏��mE�ds�4�Ip�_��E������1���@x�w� ~���D@�[*IoƺX��P�[�	��f�o����Vyo�7�SKH��~.Ȣ�K%����w�-0���Ė��i�s����9.�|�͋����+5^��AB�������Y�~�H��>�u�.(��׻1��M�޺�)�M�{���X'�#�U�иl����$Bl-E�*+61 D�_��K��e���ib��%8��c�}>�>����EbV*�9N�9R�.
 gwOr]� u��\�I�B�PoV��٘��m�l����E2�"بB�]R�O#i�����T�s�����p�P�Q ��t�D�]�M'����9�*c ����6%�t0�8>	 ���uY�����R8.��DX��Ҋ�����=�D�x%�M���,Ƌ+�g�bX9�	��n��ٔ�uwq�a5�/It~�Y�.�u�>�_���-t�t�Y����q����RT�E���7���sS��I%�J�-�x.���Ё��3�4��}�a�e�8��zo`ڊ���}3�B��!�<�-FK�(?-G@\��⋑�#&�AƈJ�O[��^����������w�7�˫�� K#-���r�
�-Q��׳�k�t�E���?mX3�Rɯ��"G���k��r���9g�emV�b�o>ٽD%��8*�'�E9Myv�,\���r.��e��dhD2?�Y���z�oԲ%�
�(F�b��B=�6���3�S�?�Zi�"VMM%�횏YS`X�]�ܜk��,*�����W�ƽl�݋�����:�wO� Y�9��g��g^�/̶� a�����N��>��9vQe�U�1� R���,v	��r��Kd?�E��\{�����T
�e�MhL��nXH��)B�f��2�'������/a�� ,� �[���F��˙v�u
�X@��޿��?U�U6��.����q-�P�ԫ�Y��� ;)eT=�Q��Q �L�X�����w]gv�!6�
�@뭪� E�9f*"����G?�/��Si�=�����vR�11��:ţ�
�}����DG'T��dZ����EX�%E��&��|ʳ�>遏 �̼���M/D
qy�6:���I��pp�q�8ٌ��u�8w礐J��#���ގ���Y ��ܡa��>�35x�B4�L��,v\�p���@\�`�>p�-ȑXcF�E��y�43M��6��3r*�q�]�n��{�k�<�#��V�qW��?ա@oz�{�K
E&[�
!�tCi�Mޅ�,�ד���F��{�UU���9��Sq�X�y�~�\�'�:(I�V�d-G8�HƙeY��d����=L�� �es���佬��c
#���ǳ�,�h�ļvU��D)�#�9�/;T��T����8&��A�Xy�׉��=���ϼ�6�1X>o΃E���B�(@p�5�I5��h��lg��S;fo^?m�me9���%"x�`y�l=��������xd���AZ� �>��)_�{?�U��0B��Z�?�7��:����4�� ���>$����޾\�X�^?md\� |��:���DR�����7;�_�L��3�Y_�V���/��W�N��� �߷��4�U�����o���b��q�/���Z��ls��adaS0��M4���%��G6<' ��:�]~Q_f'��#���]���7��m���|��h�y����\}�;��y�<a� ;���
�T%3ЈC`=V�
)KD;7���XD;�Ɲ���V��Ķ{�\��	�$%ؿ|M�G��D���z/����+�ӫ����,���
�e!"�$�X!õ'��<2 �s1���@p����$�'W/��t�/���v�(���[�`Д�v���c���sC��G�54�}
'�á�����q�M�ϻtt�
c�����9�*��QU�XR�%�Ueq�c�"}CIe�o�xN�����g"�1�&'8��\���+������N@	�\��Mx���Q���.�} ��Xc-��f�,��_K����r^�W�9��B��ϯ3Q8n��-��FⅨ�ȣ��k�~�-̌?����� R!:P���6H���^��ɦ@�N[��l�}I�7w �rSi��yKA`����?����?u�7�Mx���