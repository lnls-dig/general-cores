XlxV64EB    14c8     800Q[5���4V\�Ky+����
4Y������&�w�5�6k\*W�B�#�¹ "���W�T���+�]�M�?tS5#g����S���Bx�|��a�*���\�$����B(���Qj�/8���G�����'g��]XP���KJ��q��� 9z��?D�b)�M��K�M�.�Z��t�\�V�Ze/���I��m+���k�i��F<�#�t�K��N�e`�CU)7���ג�^�Q����_�
�j�
��)��Ǡ"�vƇ8�j�'=c����%������X�'�Y�NְN�g�~5�������m*�~�	Ѣ���z�k��S*~%�I�W���B]QS���'>�"Z�W�6�9�B�4��=aC�p�<DRM,�VJ)"�ׁ��&n�dVf�Ԏ1l}�N%�O�$i�"6$Ҧo�(#\��y���ϛ�|�B��,q�zj�g3O<�,��)�;�N{dذ�c���r:Y\$$���&1}���r�}@_�6����H�)�m���	�ϸu6��=���]=pg�'��2�A��P��4�H�{V+{�=�$=B�3s֬�zm�k�������bq����0���A�������ǵ�:��л�b�	��03~�֫��M�y��2X�����P������EIڔ=3Q�~(8��-FG/#׸T4=l羽�
6ۇ����Ta�u���
�dT�9Q��h�\0�0�h��yZj3Iٓ�Я��������"Eh�P��D�[�4\�4.,��{Vçm�e�>����M�p��������j�i���u�1>�p.5T^0*5$Qyh��	�^k��� X�.�t�"v���Y�|W3&'eC�+�q@Df�哧���o|�����P@*�\zz�˞tHS�4�ۤ�`��ux�f�@"�>=奔K~��}���cp.�t
+��H	���"�I�p��޿P�*��QBg;�
�á�W*�LH���/���?�k�ˌł��;?��"���U66�H�T���֌A�[$�-�!���l*������rSz�I1���B�JH�-S��y� �%��Q��B�.]�+�tzț+Ϥֳ}���p�[���eR��~*�x��w�|h�9������p·��k8D����E�����@�L�)�E�Aﾁ
f���*)E�6D1qz׈��lq������.�v�kh���"L���8qp��i��j8�e|
�ō��������@���PD�+�t��f�C;?E?6^�� �&��de|Fӌ���f�rQ�I�$Ȗ�{"&�	I���w�v�	��V�{�-�ܛe��YƄ�J(!��i=��I�De��f�l�����~��E��4��@�^2E�,l�􄦛�LH�R�r��.��tٸ�w���t �ѰiԘ�Lo�&���S􊑓0���.g�Σ���Y�(ǻ�m�U�i8��kqճ��Iz6N�
C�x��Y|ɱ��&w��{C�U7a��w���˾���tB�V�[��X�cڠ�U1�6pd�Ʒ3	�	)`8����%>^=��ov����Yo/m�-��E��;�&a��Q���	��"�=��R������7_ɑ�o�6���qۙ*5Y�L���C*ߺ��B���K�Ba�Q| ��6V���z%cxK� >���a�;��I_Ǜ�@6����Ə>Y��W�ѻaE>�K�tE��@�º��A�O�X 0�R3#;�2��abl]�qK��	�1sI�>�^6z�-YH�#��W�Vw��ȼK�	��������`"��&�'J�#�IEU�
�ؖއC.)D�|l�֪Ǿ����D��k=p��b��@.�]�
�hvv��T	y%��;�@;��+�c:�� �yBs	a�>4�z�����xʛ!��k�Q�E�덢����hi�{I�ݓ?X�h�aJ���QR�����Ҕ�+�ܑ�1Ǉ ۽2ş�-����˥���w�8���%�Dj�������@&S��c���c"}-�y���K��E�%	F�ýNML.�O,Q'