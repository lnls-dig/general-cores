XlxV64EB    9c50    1610�z��+��Ŧ�>�����vs�0b�LŖ��y�䆖���X�~mȝ�+#+w�C���Y�J��4�ք'�C��h�TB�n�P.æ�MN�Y�4J�q���M�dgJ��R�38YnEܼc�|������?��I=����t���+ �'x��-��$�F�����?�h��ͱ��:���ˁ}q��za����<�P��/d3%���o�t"A&J�a�$X׻�W�iOC�RU����'F�p�U�~�Ʊبd`R!%�~�1?���070�">�� �&�jK��}y ��Yﯧ�xH�qɥ5?t8��`��ix8]��EYvH�J}��N�;�a�]N���N�3rl��؈�S:#z��P-��ZR�`^��D���ǔ��"�t�
AwW�i��K(a��n�b��t:bo|��[}֪6�43
�7�U���ۯ�Hm�W��Z��]�ZhF�x�"_�U���?��CM�<o���\��z����	VIPB-����F���Mv7�w.����~{]]
@sD�(���jq�4�x8V�\���Q>����ڈA���y��� ����.}yzA���eY���vZ?�H�5&�!.�$�he��Mʟ��~��F��<QXF7mp`����P֥��j�_���˖�����%G�\�O��=�8�$��Oȳ����|�B|뗲�R��a��6�h����2�%�f��E3��=���T���mʖ%�=RJf"?�AY�4�F��>x�v!�SR��� �k��E�JE˙n�m��C}��(��J>Sr���`.a�HHŒ�-���Vخ���68��e���f8n.�]N�)�^UV�fsg�������9"l69��Z�tl߄E�s��u��6)\��X>��^�R�'O8�ꢽg�y�ZթY��u�=�(����dnZ5�
T?Swu���e�-&��n�Nx|�S�5c>Ǌ�ݒG!e�e�Un�>�Tƍ�R�� \HsZ�t>���#MN����g'�� q�w�4Y]��k�2�1�/tV�/R�?�ty��I�4���g9|��q	�b�M�퐦��d���")�V�� Աܝ�F�@J�Pk���۶

D`��W?Pjs^�U�����q'đ2/��>��k)�h� ��l�|��UˬT�K�c���+�-��g
������恒���<������1�;y*��'V��Bvޛ6I�w��l�w����:�G�@�����u���FH���Kb�n�$Н}F�s��;�|,6)�8#�_�)�b��7��rA4y&+ùF�˜aֹ��i7Y���"���O��� �8��:�.��q� ��2�~ۛvXb�ԃ�}E@�؋cu�Ż�y���$����[����� �͝�p ]��)˦;п�
�%�Ƴ�3
m\|��tW�y&�{"ną��������2�c�H,4ww�va� Ff��@�5mo�ޱA��_�UvjS�G&a��Ð[������ޚ�L��!�^֣�,'���F�|>]><�cy���Ѵ�]D��d�B�/>=�c���!B�K�a�����;�A����9>�.�t6�����G���3�%\ИХ�"m�@#��;UE	cY�O��)�>�i�=e��Fo����b�E�[]��=���R�逗2|.�Nc�27��<�K��5�JHt�̱u5p�\m޿t���ZP4�;Ϋ��Yt��~�#|D������cM ����v�����8ܹͺ�QW��EO�:�e���?�W)$�A�}b��x���	�,Tsh�������\�MC�`f���;��Q��P-�,mSa���V�g����O.ȝ���AO��G��C�\@@�K�V��-♚�# /ޠŰ�]H%��������xH\��A��ƌ�2b�6��u�{S��O����YȆ����.����1�i��LX�:��Pc��t��W�ʀ��&/��]E{"��\'�[X�^��|͒@z�s<s��r�m��p}	R'�#��0tVO��u7�$��7v�U���&�ڤ��H�B��$��^8����Z^Ox�Օ��j�S��q]�$9�F4$�t����G�
��a'O���9�5�:�����d�#=��`�1	
j~d���:�o
s���z����ZM�2��&����%;b�� ?�]?^%��PJ�G�`�k� �H���D��1D�wz�KMǤ=VD@��n��ށ�݌��Չ��5�h�B���+q�?����H�k���Juȩ�a���ɷ���AN4�S-�J��l*�8�RtrM��Kd��(6?��!l����d����UZ�oP��`��\�ח#x���KP� �@�M&����@
M7U�\	̲�������-�ǽ�L���"��2��g�=ULd�����C{#3Y-��H��a�=DGv�>�K��UBh7K6#~ÌP��.m^P���^M���3��x��o2�Z�����=�5=��G�Ku؄.�da�d�{����r�O�?�O����H�S[��e���I�-f��kZ�
x9Q68��3��l&��6H"n*��𞨦��5���g���U�T���)�#1��^B�/�v\��������*�E�;+S��!&�ʐ������T7���Ij)��Y㜣��1"feHS ��:L������� \�d��c���g��F	�J}��!��	�a���ϭ&�ᨋI�S>���]����=޺	��\fo�F�Y;���H�[�/
��7�Q��O�uq��EZ����Ӻ��׸G������2�; ���wt(���rBg1� �O5����(0�JT���y�ľ��zw�9�u��hI̡�Q��#s;[���[����"Nr�YwJUۉ��	�/f�(,��uM�Jsj���k�v��bI�Y�WO_Dr�|1�XP� �s�~��l6x�5SdXm�w7��`����|�	T�T���T9���YlQt��~�LN�S-Z�:�-^6%�´o�ߦ~�z������kJ�dxa���ǕI�&�*jkK֓hlg�l�Q���xY;�"f�����:,������_��;>�s#�%�>�[�s�T�L�����9�bBO
Ġ&�`6U���������U��k��,��Fa� ������{�7_`ϤDV��We�'��� ���~EN2��䮾��?#�J�-�x��P���#�-I��>/��_��t��c��rs���P��� ��I��̙� `���2"��K�Kϕ�y%w�;\�)~�~��~�|�V˘�#	�_�؅s����\'��?zW��a�EZ���$����1X�z�Du5�]/K4Pu�ntc+S�����/MD�z3<��^��Ɵm���A[���4*ӌ���i��������a����!4l̠B��N֕˧��\}tiIXW
���B�9��q�.z�^�ة��ԣ�8F�: L���{����#���w	ª �0��sg�����C���V�}��N�����t����C�(��0	����y?�k�2+ό�j��d�,?����BK�@� s*61�vb�e�`�[��v�|d�_�C\I}�w%u~Q)���x���q�R٠���3�A��Ȍ�o7�@FRmx+�b�V��7� /iN^�����b��)UjE��`�i|��ȅf�C�_W~�l\�hiu�T�=�E�ş��Z�(˒>��^#6��_Gq�d5�
�.�����1"=,��y4� �w�׊,է�V�P�J�Y�3���e���q��B�d�������C3�� `
Ī��"_l�)u���Ȧ��G����JNOKG�>�^�����h�����-~6��R.�w�OT[��Ū�!��ؘW�M0�rC�7��O�ʡ��~��Rou�=�8���[��7�9V�CE�T��Qp����Y�Ժ�s�Z
yY\�������Ou�sXH	�i1U��G���鱊�dހ\��VoO�3���4r�?��*��ݜ"F蚰,mkfG��U��9ʥ���0Y`�R���xۜr���^5��i�xo��b=� ��\�Ê�����֞�d��v�wЊM#U�f6lA̅�HǞI�|6�p�+`���7�8>i1�~������)]q�Pk �QEmb�U�,@���n��JQ�MR_�W��J��ܱ���4�؏�$2,�(B���D�L�yV\km���`��kդ��ժW�v��b/17a��H���z�ʱ��z�����^j�j-14���.����J�5ĕ�;wm:@�veDV+�b?׼H!PnS3D�6ۢ�A�X�oU��p��w<���|�8ol�� �\s�@�-N��o
��E�u�U�;K�Lu���]q�ż(���se@k�~��թ����� @+�e�D���
�+��>�>4:7@����'��%!���Z�h�z����j7t3�=rN�'�e0?��%�C�pe�@�WH��8q�u�J+���n1=�,�ݶ{��T�_0���4����O��67g��M�;��Z��>b:�^��V5c����	u�y@c�S���*�.Ud��q.�[�k	ES3U�z1��{����g��-:��$�x�8s8F]��<3�����"�@���c�-�w Et�VJ�˚�jW���x�X�]X+�I��̾�_�%]Q��Sg�X$���M�<��W��6���������PV�ZTl�8���R��\�l1:u�{2m++}븂<xi$���f���X.^0F�H�0��=���[n�d�o�Vy�a�Qڡ�Α]�預�Ӕ%{�* �TQ���K�������Sz�8�<��c%�(e�`]�ϳ�I-�Dr��C��>�;�Ҩ�M�~i�{���.�_t��zŸfp�-�0��O�'��X���j�=�u8����^���hj]�0�}G~B�O\D�N��1@��h����r�9U2��H	xe���[Nbp��Qo��#_=M�k�ԓ1i�cOŖ8	}p�nc�� �_��������d�+&�v�m,�64{�^fB��>V�&���9A����
�����p��
��V�0�l��)ȶ=�ě���'�1\��+���#��A�,�
�t�y�|�[G&��c�-<,��!.LIre���&2P�/ʤq�i�ؙp���R�i`YzG+�K�:��H8�94�2jH_�w��d[��s��b������	7V0p�g^���.}"��n�X7.�ZI4�b{2�na�.�+�p�B/#��ػ�%���C �Hm�#��D��:&���§�{}#��X���u��.p���Ny��\R�X�D�f����i���J)��{�P����0��9�i�W%�\J��m5�~���i m;&�u��_�g�f{��W�.3����ێ���%΁�Q��t�_~��G��$ߧy����˪}��l��S
tj�k���ȏ<�D��6Ϝb�ݩ6+0�mt�ͳ2hr�u��q(Җ2�æ��H��}v����$Vu��m��o���w�YZM� �3UJ����B�;�I=%꺎Z�v�%�s����;�zۚ��.w�