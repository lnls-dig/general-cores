XlxV64EB    8fde    1db0��!xlb/�=9�#� ����kb�X������S�hž��U>�$�F2�;8\��>��ځ��G?�Q�u��G|�tTnIܣ׹��9�3�b��[�	$Dc��e����<ƙ�/p�BKF]�����$ž��Μ��(��굴�k�0�)��5�AQ�Λ�&���Ptm��!3$��s|W�n����6�sz�fv˒�xuy-2ˉ�L1�i�p����h�Vn!+� �j�f���*s\��1`k�I~�e��
a���do�\�b�p��q@4������=���3�G3��G��(B���V�=����¸����j�*����$�[:Ѿ�&ޕ^�=�����r��G�Ci��B�o-*�D&�F�&���� ǯ~ȩ\?��%���4�p����vN���r8�^��.�wbh�#]�-�ZE�w��<��ٸ��I�AU�z�5��v�s�)��_��6�@��ʐ�`B����Xh<Rcݴ��@��':��-vw[0_#�k��d8�MV]�؀f�2r`��h9��F:��Bn���9�c_+��v']J=i9'�&�%�qp� �+���� ��i<�8rBbO=�3*��1H����z�hT�aBDH��������lg�?qJ���jY�Ī��r�2���(
�6ˏ�e~)��㳍e��e�U��1\>0OYD�Ѐ��):�z
=�q?g"�U8[�'��Bj�B�ޣN ��#V	�V����/_�c�>��� :~��$(��#��n��M��=9HH��馿�=��;>�p�4��k�
!J�m
(<��Ȧ��ϒ+�rl��S9�Yȉ�9El��x=���j³��#��Pp����=z3z(̀�\|���5�8��l��D��ӣz{+�Ǐ׻~�#���DQ�̈��_���}%���<hB�%��JJ���X}_���F���A�G���]���n����M�[�r�&_�k%�]da���+Ō�P�+͂Sg-�]����T.B���Y�V wow�j9Qթ�LB��)�I��Q�	���϶~+>m������������l�|פ#��E�mUQ˺ڬ:���]ǖZz��Rv�]cQ�I�H�����o�{���j�O�0 W�]r)y�d�
HPm���Zz�n�nY�����F��u*IY���*�F�O�Q�h^��lXq/%��B��*��v�0,
Q|�W�ML)��T�
�A�\�����B8�/��ˉ�M8����\�V�� +������4k�G����4��\rd��ޗ��Qcg�ㆺ6�|��䲵K�!
Er�w�2�8!��1L������K����Eu����F��ނ'D���\IKר!�Z7�af?F)й��TJ���f<�U�o�H2���j����'��I_�(UtyL�� �4e$q<|������5f��ʄ���K���s�M
	���#b��ϝ+x�_^�c��2�8_FQQ��Ki1q^�u�
{�N����)̀����E�PT�^/���e�&P�P���j::`c��k��@eɴL��!',�-Zx�h�u~�F�����;rp��}��H֚�5�V�,��ZW�V�y��A��+F�Ԙo'� ����O��%��[ea�u�'�����ӥ��O�r���/���e$."[��]B��pƔ=F�l�b��h>��L�#�p3��E��"�^yFP�lX���#~�`ൡ�j/Ŭ����:�wܑ噁!*�H�\�	�citߕ��P�7�/B � =Ɏ��d	y�퍫�!S�r����&mkZ_�<��N��BF����p;gm9jxǅNIRV������aW7c˰Zܺ�П���wpn��.���|�QI�BYN�*١>Q��p�ʱ#I�'G�T������[0��_T[�P�W�6�E��es���A�epج�'�m��f���U]�S�7���惩���#��Q�%�x�k���r�fC���t���D��	\�-��':u�3��b�-��s��^�f_h4��^V�=	�H�UO��`�6h�����N�G��r</����o L����+��XH?c���ce˶���_����2�����b�AD�'�5XD1��
$T]㘬�;��}<fJ�"��0]�5L*�ėԣ�rV�Kvirljz�IC�_��(���$��h {�O�j鋛V����n �
%'.1��|�#�����!g���
�-D�Q&~C���[�\*Ee�MC��x@sn��R��u�O�," ���+ܒ����XO�c���1/������L����;i�.�e���o,�9����w}&'6�cNx������Z>Ê(��=�+�ƌ7������0��|�7��H�_�x��h�L�X�6z��Ͳ<��Fdy��/&���~�ڢP[蹂$�P���)�g�̱�.dt?	3�-#������P�Q;���g/$��e��!:X\�v.�dշI��ϛ����t��me����]�3�t�qp�h��o�or	{���7�`6:��T�E ����ͭ��o���(5�c=VdN�i�!�ˇU���[7�h6�1�^��N��@3,��;{V�(��wY�)������f��ź�Y��F����>��NZ�b�4�����_Bbi�TqD\�r�	����1��O?�@�]�
1_�d�^�6Ê��\Ү�i�������>�]n�
��5W�$
0�^��Њ����I�@Ƴ_�6A��m�2.���O��"8')��~��o:6O�J������ș4�.g7r�<�2�P���]҉A쯳:?;��縏���B��ݜ�L��0i�s�k=8��t��x��b���S�$��x�K�/��Đ��%zQ�J�/K��=Րɫ�ғ�X�,�;�`E>a�4HD��%��k�]���Z�bԩ��V��,�A�B6�2	zi���&�VZ�@� Ŗ}�d-�"/�P�R��-]/=������Q��t7F���i#��a��'_��t�	�����ち��<�+w���z��W���YT�a~�_���Ah.���)cG�&��v`��r1D�{ju�S�8�i�`l^�YɔB��`;��ЁF�N���w��ޛ��x��Y���G	�u���uӧ���d�o2����T���S�ͤ~���!.��-ق�)�\̆�V����#F�� �$�ZC��g�1�� �8�C�Ӈ2}-W��i$(=������WVF�{�.���.|�{:ҎR���\H���o-_ep����@�%�_1,r|�����#���2��˘۰:���[�E�lz������::�lz�yZ�����ʙ�O�����-`�:���q��kv+p_%�7t�������0�����@z�*P\�jtA�4á�rA
x���0
��[���4w�!��BV��`�"�ܟ���{��~�U)�d��J�&ǒ>I�V�)\&�A^�LިzT����\��I��8h���9N�������+K:��+�'��n���9͋��^n[��"�&��|v���sP�m���6$K��̩^$�a����q*Z-pa�<F��oN`,|����?!0��ܼ����B����?����-\A�e��h�(�z?����k�l	�A����f�Z������~rS�V�D��Q�%H���"�d��h�������&�9h%O��?��H
i�٢��:�s��_g�/�a[�CK����ފwun��M`h����X�(dZ��N93��I���.L�v��V�}JĞ�PU�Ycq��KH;=^8��i{��MYZ����o��Vk�E���dZ��09�bu	;
�,�i��j"�B��\b��$'���2{�}�,�HX�<dһ����] ���<ьS�=���/��|�ۨWͣ\�����(�ͮR�%xt��Y��)��f�4�֫^�W!x������*�s �G����rju��-FJ��D��~����\4��-��#�J�*�R­~ec��nۣ�V�>�.��\��Ӧ�6��.!��|�Ҧ6���+EQ(Hr�e���{��������f���2��ZF�JH�q���!�����߇nց��i��Ew>�����GH�N򄷯=O@W��Z'��Ҏ�a٤�>)�#cc+��Z
�������;�]�b�~�: k��=�j��@m�O?r������5�5�'D��m�a�0C�OWϤ�X(����X�kp�"k��k�u�C�����<�\�3r���QD/�������5���kED��v���?BP���K<�(�)��l��B�Kp�Q��O.PKaX-�� e��pHb�xO��Қ)~�~?�dy'�I?Aa�l'8�A;��ئ�2̄���� !�0���В�ɮߦ�S�&�'��k�d��So���3YF	����~qy/j|�jC�y�Ñ�)���?��~8�KJ�\`����s�|Dc,�TŔL�
yyb���~�*jm2����h�X�ZwT��J{�@X���]*�[̭�f 3�7A�l:Ci�ϩQ������t�kj��f��Hp�"[�TM`��Z���Q2��
����g<h�IU�S��&`$�����G�i��=�V>V-���������_m��w
�����D��V����S�NY�bZ1���r�~Dչ����.^�Ʀ�=�b��+���@Z���<�`�"��2���6��;~�tn�ٹ篑�zxnd6�S��OD�`�~pw��\�x�L���x���V��	��[>�CQ�uE����ym��d=}`�S8�V��I3𮿌�d�B�&����{�P�^��r��D�;��~�`vޓ�}"�&��8
;�!�Z{��?��Lc�ss�'��!�[����R��q]����^����� ��3ܗ�D��Y#�	�"|�I��D�ȍ?�
B7�:�r�j6�����E��.&�kRg���Y+20߱�Ҩ��ar��#�y���lWK6���V���7Q����;�5c	�B������Ř�ji�l�~:���U[э7K>TnǴH�@(V1���Z�����%h��]����dD�kd� q�Xt�-Z��2��=2�����YǺ����N��&�	����G%�t6'W=�T�IK���]R,����-8�fڝB�C�)���gb��fa�C9$��J�JK/�-TZ�� ЙkOͯ��HX�5��]l,���d����G�ƈ�JlzG�s�.jbj`m�i�r
-5�f�K�9����Ple����M6���P�+r
�i�2k_�FE�NÆ�$�|���f9�fHcc}�W
3��+��e;N%h�#�(��,AԶy���/�+�v)��P^O��n�"B�23���ڋ��R�5�9�EF Y�]\'��vf�J�#S��<�p!�%\%;�Eo�ϰ��*%˩��y��&[s{�`ğ�]�B>JP�J-_{A���a���A����=�����sQa���-30,5�y�*�Q�XY�ù�A=n 6RB�ִ� �� �{/6^Ax2tr�z���a��%��;�w�����rkT�*��������'E3��JE��~A���~�A���*cJ��.P����m&o�̀�M�
F�:��dv�;�R��jQ���S��U^ �ы!;T��],�$g[*~����%�|}8.�
��vK����)��
}�g	���9���d����l³��LB�.-Wۙ��	�����g�EX�0E&+�>������i��\�.����`���3-�*D�IH-E�X��p�� Ѱ��ŝ���S`N���X&���������n�9	�o�M�x�*[m�	k5I����i>˕L%�ŋ�>�M�z���-�Va�Qpl���{�?�L
�'�����i��(w�w-��Q�;��9��EGN��?r�%��Q��@M�4�pn��o��B�=�ѺG�{;Zx`�sh̝��ɧ1�Y���T�E2���i�X�����A[Y�����oD.��*�ն�� �𠏵�����r��oE:1�͔������`d��NT���nD]��1�@$\PܺT W\�#�UѲ,.t{�y"5��{+EbG�{��I�V�B����O"�+m'�G��t'w0<���m@m�0��WFa�d� �#@ok��93Pr�P��7���㨟�/��i��YZ�P����D� �:+�"�RYR9x5�v)�}��Ҿg9�)��8�G�K�<��9	�h����˜�I�(����t�fF�P�7m玪�mF�j�ó�s
f<�G����7Qe�c��M$_�[TV�:����cڠ���I��`���t">/P���0G��[?:LI�1M�e|��V�^y��[{���I�p��M��B�3<w�蜥F9���6�~$�Md o#S�5U�� ����ˌn�Xn.-!����c���g3�B4�2�f���O!��8�]`�Ko����'(��߇����׌&O�y��61��/�؋ł�G�OM��n�<߱tzS{|Pc�׶*�Onr��bV���p�3zW��ד�zV�E�z�w)�t@Sj�9 ?m��꒔�)�᧫L�H�[Tuyq�ǠS�)AG�����f�w�kG��͐�F�8�yr.���Ƶ����qŷ��e�6�~�������~=�J3�n( f����(�O�{	����v��t�-z^��|��lهeP�������~&�� �x�"�i)p��2H&,"w� A���౐/����j���/{��F ���"��zg8/�)'�U����0�b�����܇/:�bd߉������D^�sU����6�FA�_�5,=���Ṯ5�Q`��g�������j��[��5��h���Q�2�a�zR2��:-YW6:�Mǐ&.����q��I�D�	��H��M$dȑ~��7���QD�{&��K6��J=�+�ɐg�+�W��=n�<Z&�p���K��F𯚩�K�Y������B�a�DJPG��tZC+��_���/3�v�`�n	��q͵�R���+t^�n<��I�Qt����]d$����)+$	J��c������P��Np0��6��B�4y���wGV���i�v��R|^�꺝��m�,��A��ns�D��ꠝ�c�g@b�b� �B��!�桃mR�e�lR�8��v���^��JW�͓�k�*���
k�,��GP�������T����7��Cy {;t�l�:����'��V��}�C�`mC۟�ʧ+�F�CK$R���(����I��n������p�!1�8�҂�rv{��>��21��Z���|)ILVL��}�E%_�A&��_�Akm� ,x9����Z R�� �9:�ز>�[F��������Cc'�
���~��lk���0��������F�L�3���Lb�������r�<���`H���Co���ﱄ��:�5˛S�#�JЊ��rKҦx