XlxV64EB    38c0     b60��6I��f�o�{q�$�I1�C%G��^ĕ��%�s�]AS� /tX�����]�%Xs횿����Aw��p��L����YWj������O$�slYf�:WR�6N3V�k=��HWM��� ��u�y�x��� ��J�!X�2%X���*�����q+HB'm@1��<���/ldl���>1��u��;�x�'v�r�qb�HJu�ғ���,�����P�UW�D���C��DK��p8��_0/o�Ǹ�S[&ww��s������6�ƷB�"�ν�W�qp�1,��O���ݑ�g!�HQU胝?�xtY/�gׄ�=�]j#L+�Kt᧫3��M,����{��s��#V���j���Q�
eO��]�`���B4_���eg�p�=/��KLid�[���
��zJ 6,7!*�GL�n^���=�d���h������&�V2�L-<r~GJ�q�2�=�4K%��0� ϼ��T��T�cٴ�����ٸm�{Tm�� �T��%B�Iֳ�}�`>Dj��E�3��ƴ<J�d���Z��n
���L���Ǘ�^�-Գ� �DҚ��dJ�h~�������E�s"�/S}��tRu�M�S�.�`c*%!ǘ�F�BE"�ix�.�:sܑ�������`��KF����8�rM�H�n;>�'��^7ͤ�
��{�����+�M�5x���B���s�~�ʶy�Eqب�(yL�]�{���K`&�/3��%�����l�	6�=�,��0�3��`45߃\ʓ�����~f����K�3i�ũ@�1ښ1�?��HY�>i�B��[b�,g�iB�*����?�{�$2�#sː.d���g����<�}FF܉n�.�r�Xq����I�{��-����g���Q26��E�=i�����6�ևߕ�W��nK�s:���&sꈆ>LUN���xh�N��N�X%���+��VB�b�:IL{��Q~��Ve*�`��ө"�_�J��������bi�xso�a�����z�xzs������n̳�@��u��U�r��xUc�x���b �b=r��D$c'BޞK�)-���ch����SKia��41�Σ[MF/3�?�:������x�O��`��w3�t>���I؍��*��5I����5`��#�g��̂������GbO�}U���e5hMO͇�^�(Q.bQ׬�b��w�������N#�]�������&�����<>#+��S��%+;� 7�&3V�&Z��e+,��V��rጦ^���R(Mt�Cw�͑�P%AȌ���H�&�������k��&:i���\���r�6q��r���R� {�C}�=��F��[ ۦ�l��rIu��E��bo͆^�kz:��RO��@KX��ؾ�x����n �4��<<L�+��Ɯ	��X�S�{�_☎r�;����-��蜲6t��n�=v���Q�� �ߜ͟&kW�)G{��qX�RD��%����5��ξ��߶���qH�6G2՛kM�į[��:���<p�t�m�\�WO`�Q�1��ꝍ�8�}����[��ˇ$¹�4פ�^��'@T�afT��b���%{36�X��߁>�������$�0��Ƈ�v�������[��W.�^�a4r��<��UZggyt3֩3e4�a}�ڍt��"��_�h�"�:����i�I��j����BޔS���S����Ƣz��V��E'@�]��`f��TzI���;�n���f��Y�ox�b+�Vc���kgZŀ탃���`��x�`��a�b�Zb�o#ZS��:e��.+4���P�:��d���x̶�X�5Au�f$s�Ғ���)��R�sB�r�cg�L1�ҵ-2��k����4��#�e�~4g�0�'��k�;˔�m�t������3�����;��z��R�,����q8����`az����a.þ����>�:�`�Nl�gRڒ7�Q׉l�#cG�At�Hi�$a$2{eC&�N�pQ����,�cCw��c�հ�`�r��7�"���9�$>	9��x��3?/}����K]Vv-e��zl;C���v��HY�j�w}�9#0��!lJ��r�q4h���ѩm�F2t�t�'�o=�D=�o95�=��"H��o�(	Z�阚|1�r�L���N����c�!������I���S�0�V��H/�� �p�e�.�-*Xx����݋H#��$"�L���L5�u@ѹ�[���+E�٣�7��@@��ed���J2C&�<�İi��*d0���Ɯ=f����߯�̉�鲫���2�!�~G[���Dk�j����.P��a3�;߬��e�\�k�f��ܙ�},2E��!�PD�%X?د�U�؝8$Qٴ�� Z�vY9pZ��wA%�,�@h��o��c��Br�!�ä���ػw�h.���P���A�d!�wK#�
��������ɿw6�v׫v9�z��a"9a]�~nL��atq�F���aZ`"����n/����bB����0�`
9	_�Z� �����:�E"��釄+�$G砝@to��AWHo����%r��`�f<� ����} ߴp��'Uz!�BQ��]���[����k�%b�-4a}Ԝ��I�
}�fBq��b�����sF�3���� ��酇�]��f���_�&�A����qrHK�S��ƨ �*,>��+���Aa�qa+�3}��'��ӣ���M���T��4���0���	�c�z��k������|��LN"Qp�9e�)�IAR��oS_CmrY1�& !,�}UO��.��g.��%L����3�
'�