XlxV64EB    fa00    28d0
���f�6�=�:�d8)��X���H%/i�iPx0�`n�������p��τC�\����F���B_�8'<5��t���lv����4VP��*����r�e��������D/C�j_�3��ѝ�����"��4�����a�1B��@�� R;��hX���?��q���|x���R3b>�'�T3�ۻzobWڮȠ��z���
NZ5�6�57v,r� ǱY��{,�f�؃�=�>^fx^�L��E-��`�`�PJ@9,Ν#b�KO�e��T��ao����)�8�+=~]��-Y>�ʙ���k(�ב�ڠ�4�IS;�^Է�+J�t~������bK]6� �>Mj[��k��Y֞���6����1COL��g�U��>x%[)��KL}�B(}4jyr�՘�(Jo@˙F�GN���V��k;`J��Q!�44�K�ՉV-FMں�3��ͨO�Ź��X�9�&�~K���
��AFr��m���5��T�R��-x��0�MLF�A������ N{�Zh�'+n���Ҋ;�����V��Ӿ�A��	������I�׷h@�I6�oԆ_y���̰�^�bh��	��)Ûs>(��E&M���5KȬ賭 ܿ7t}(��-�(��Y�b�(M6˛
��*����ϹWk�}�X~���+W76~e!:�z68?�N6��K��7��qh��:�ޭ\�,ԉ���~F �m���F�([��0�v�8�Ę���N��q�D�K���	��H+�kL������q�v�%Y'��V.�
-^S�Is�0$���ٽ{��q���Z�7ݵ�L+Y�k&����%}N����ٖ̍�Y�2U�Y0ܟO�v��"�a�/ʅ]t�M��Ñ��=@�?��nܩ��b๲a.��2��9Gۏ6�H��x@��C5��D*����퓯���e���CP�@N�#�wjx�
���=��UC���:�ua ������|�r�-�����/H����+�hE[.G����q���^!�u���o�����q5|Xa�Y�
��1�+r��\/H��)5��]��7Ibյ�;��>j���.�0l�kX�DM���G�4([ ���ʧ��.a�W.���5i�����WI�?�fy;:���a��t����J��6Z b��#۴᫃���1�q7�@��V�s
�_:� (�\:HAu���f{T�N�݊K�m�����fv\�|+��W86�af�����T�ø���ځ�9�
�=��y�����w�����L_�Q�f�!$��+P�L>//SV�U�AW�pǲ�r�P�����w8��?a�����2���G3A�ԉ�w��d���Q�>l|�v��`!��R��Љ�-'���T\#n΢����@*m��,	%IRd����6,��Ԋ�c��o��f��"��fJ+��%�ǘ���)5 ���<��d�Ñc�5�'�0���>c|wvlu�DN����,R�y�(�u�����\�xȰ�U�0 �SA�_S��)'�d}�#׏6CI�NqESt�22��$��.s{��u��4�	��(�l?ȹ[���;P.xF�+j��$G�7O��© Zk�V4�|�H��1����L9��\������p�q�Ri�e��>�;�-2jxg*����/e�"A�r�Ҭи@�%���9�c|J��:6 ���,���7@���U+��A}()[Ba'�
�oO���{ʌU��"yE��n���wOŭٜsq}���(7�ތ�0_/2��:E���c�g;��j��8cS��N<U�B06d@:=�%0ۋ)�c+wy�G�	��M��^����m��	�m�a�yIp�@b#B��-K�$�9��*px� 8E�Hhw������ϕ_�8yu�Q3@ˢ��炣b 6�fd��c����B1+�9M�<͇�T���)��J�	�z�jC}�	Q��2l#�:���Dc8!"� S���[L1y�ۑ�n44�U�4u]R�r�-4����cq��Q��a��I����P����][|B�N�9�\�N�_�Z0��V�Wt�[inB��F�c�r��U�T��/���NbL��)p�Y�n�Lu�$Rt�C�N�6�����9Z�L�rp.�#7�K\�8y��i1�/��\j�bPW���۵P8�s��Y*�7�7��\�UDH��Q7�π��B$��	s˃Y��z�Q��T��wi�����d�ckf�~�(B`�v��3�u��+���{������]���
H!��(Ө��=��0�x��l=���N�-1�\H��z8�@;$�)�D�_��~n�G�*�F���a����/���8�HY*	&
�g��A
3�trE{�w,���f�7��	9��?�2HK�ܞ���)��O��F���
^���-ky���cI�x[�($��+�n6�z���e�u�H"Ҋ��&[f�6PpBߧ�֘\I����a�ߣS_�(k"�u��������3�k����"W��m+'���[��*��/�S_�qb5��0�&y.2%�@�����Y�t�ꍉ|B�S���эX��nR�
O���'�K��i�>�XH�.Ao��w��-�7���QyXP�-/��~̉P��⩛���d�=�<��R��`ȍAY#5��Z$���Y!mFȌ�J�=��i��1����M3k9�s�^�W�	�9���(ix1�y��O��7�pū�$�\_5��EU���;�{ �FȮ�a���ЌD�@���\��\�4�J�k�1�!7�h�V�s�=�|")�l]46��9��YҞf%|(3���]}Z��D&��+����݂���T�B̷����4+I�]�fh�Z/��H�P���X�`П]ڊ�����x�t�i&_$�A���j����4p�p�փL��ţWoiUjX��7y�xw�D�x"&���-υ��NH��U%�j
�f����23�.��yz��������^`�֭m�:��\���"�W���֛��0B-ſ�<_�
���m��RxINx)JU�p>/�5���]@���%g�e�	��5�|�Ѷkh�?w�X����&���E�p:���L�s����Q�S�r"U��mu<^!A	�� ��B`"��2'����g\~���fLJ�ȩ��Knf͢�m��~��/�^�A����d��|����ͻ�՟����I�����X=���Y�~�z@�yW+x����r�h�"��"p��0���$5�.�G3�e�ar��s���7a!Ta��1�d5g����QP���7~��f��|;v�a'GiT�����q�h=ߖ��x�\!-��A��͙������Uz����XG"���C¬,���qF3�&�}_���6�����Qc�F/X雤k&va	�<���}��5`��x�V��[��ī	Vu7"��6\=@�T�P��(~־�SBK�f]<r_�/����5
V�N��V]��k�1��O0	0�Z�Я�v�A�QO�o�~��w�/鹷��b��S�e6��(/�wK���c_��9�h�[��g.���mZZ[�Ys^Ho�����	酔т" 0�4w�I�$=�����<�1�x8,DL9��^|}�0�!ݻ?�v��!�n/WW@�/�����L��zb
��(S���f�S���)�I�EW���j�*����2l��uKBĆ��2ru:�G�I=�^�U2��|Z ���s��u��xI �4�Y7��p)�Dn�C_���?oq"3�����Y�@�ޜ|ݥ����a�e�c2g+)��c��5�oS����?�����|�<J�8;�V��e8�H���\XЌA��R�t��k�7�L���ƹh8-7��߹ɒ��8�3r3�?:�$A%���}o��b`�~�F0��K4�`��Pi��di��׾z`Z.��l�C�O�m��Ƒ�u�s�Il�w_�"V<�7�>����%�ݵ~�'��4H����xVL�MeE�	��x����k�]�eN2��!i3I�Rya��)�"Mb�B%t0������p9IY��'�n�#�ލ�:�+�3����z<��0�ӱ����o�=5��?*���2���χ��ds� ��6z�;�v�1�ƽ�7u�!ԧtU�(�[䝀`&<�����O�[q���N����i��۳��#CF|�Į����p��zd3�q��/n����[ݬ�@����5�q�.�]�b��ֵ�i�4��%^��(��r�_������P�k��E�,+o�y�������%�P��ƚ�)61ז��������y�ݏ=}���ݢ�B��u`�t����o�-$念	����n3{0�W���� �n��j��E�>q�|O�����I>�Xߑ~h� ��kh�ZF����޼�g#���f�& ��֯�i���d�EZ��-O�����s$�;<��V5[ؙy�R��G��:�S���|�Zݲ��	l�$� ��.=~"K�]������%Mme��������F��b��[A�D�[��A�p�B��c������1�R�gO�wm�ǡ~�ː��tj}��KJ��2a�ƭϗL"�| ����l�2F�K���{�b(��/uH	���۹�$Q���C�9��,x5�L?c�������8|:�-�	o��0%#��i����P8<�9Yi#���HL*:��	����#H�g�+(��ј�#�����5��b��rq~�Ǧ��v��O�ΜS��,UW���77����*��4w,Ѻ��5.�?:���
�>�ۙ����9o��Q7�>2�$�����9P�W��-���)��Z�ۉ�nHF��6�]�>��rA��D�<�l츿ks)~��A2gV8z[v���2�a��A� m��ps�|��,��O�b�֏��A����ۀߪ*��0�)>)ѥ7��7�����وxQ��K�>�Dۛ�ON�2������,�0*6e��ǲh�l�d?��jncJ+A,�G�����Y�}��M-Ж�Bd�y�����\R#�u�!� ������$-�>;V_u���'�uw�.�Y��ÃM3M��A�4�2*��T��3�63��JF��,Ix��d+�~=T�`x"�3�I�@�P(-f��
a��շ���j{��֣�r!�!-Ј�G1_���A�<��F:u1����O1S3z;��d՚��$���:�J��Ks������>�{�-`0���l�_'4��H��4����[ 8g\��D��J'Eet(8���o�'�{jg-�(zÈ�䓟�� ����bG�B��z�ͤ=�q\��1�s[��o�����A-�jU�@\�!c VX ����x�3���g�a��4dm/xU�˹c���'%��W�i�T�Q7�	�Nmup���n�!-0��n��������+5��������z'=L�;l����S75>$M��=V(�����1�Ю��`A�}������Ō��7ݛ�#Z�G�f�,�S����~��(~���I5< 8܊[N��Q��$r�Z5����M�$'��F���r�OP{�'��әevX.	���<1�%�/?:�8�P�yv`v<��sJ��k�L7x�F=/j�MUTDq�[A&a�ۘrO.�����ߑ��H"��������W�A�м�����}�(��x�|ٵ�hD��8�Ćp�H�Q���k	�`�Y��B��_f�իN�;��#��`����A���S��_=����H��ꍚ�Q!�Ȓ2(A������-��3��5p����0��a�D4m�w���jEC+;[2��{��uu��&Dv��F�6J��9^V������Q��ְ _�h���K�d<���=�8���}�R��y���mzH����W�7�T�͢L��vDWr��i=�[���	� �.�ݼ�ò�$�A4E�{ѼY����E.�|z�����>�����!��"�]���VZc�To���v��m�����k�����g%fg�?��EЫ��zXm�wsϔ�@n��?��@\��X,���W����h�U/e5�bR�D�qd~��%g��3�c �T�Nn�<:|2�#��Nt�wEv	�W���:��ޜe�e��)�J��tL$��+L�f����������
�mrd��+�~�&g@pJc����1.�.v?"{�%h��g�U�}��)��q���Cn��7�RT0~��.�
̻�/C2��C7:>�k=����X�R_2�Ѡ�E��e<�,N��uxzã#-�P
i��Rβ�����\��"�Q[������.����i���.pXa':�ל���d�)��
OH���E�׼՟��a$؉3�Q�^�Y�&j��,h(�\_o$>�G���I�+nGL.$�h~`Q��_d��	>�ڮ���b��ڳ�Hl_1�k
"U�V�C��BHߡaՐ��,�;� ���fT9��|H}��r�_=:қ,M��4��{ >=�j�K�M��	�.b���"��.{r����G��&v�g�Wg�Ic�(7��Z��@����3�	��Fb�f@O�ʼLO���!y�L�Ã��AE��Z����#6�q����.A�n)gr_Rj�:���6�Ғ������S�~�
�����^nX� �6#��
�� u�C};&Y��Hc:(+C@͵�%
DS��+cHԉmB��؁�=��p�q��&�j����خ;{P����ڊ%�	f ��4,<T��\���2�,M��Q���]O�S9��7��������byjOZ�q%"���(
�"6����C�$R�	�u��R�DU���j`.N {T^[��"��{�4�[�YF���#�%��q�<Ғ��������X֜Z6V��r=1�hOT�'�C��s�36p�]�1���v�i��ث���ߔo]`����M+a���]S���~܀��"�_ ��֬��zo^%���ʾy�~B�W �*o���~�N��aǲ;����z����3p�]�]��f�h6���B7���m-Q��7�X�׬�?����;<J�ʿ��-��*��M�0��0�9=ξ>i1S%�Lɠ�E��y*��H��@�e�R����+�1}�
�k��A.�	AUt{��a%f�aY"B��WE�$�kN�7-}§9�ڂ�G�K�Qh��u��6�tA���ƹ�tG�J�m&Q�}�<�tx��B�@x�f�u"湁:cSP므R_��B��o:�B�K/��"�ܝ%�4�-P�j�n�-X��;Si;�
򶝒�܁��f|�x7;1��D�j˛l�H�4�x�~��rH��^�M/�Lu��j�%^�kg���g��++��\M+z*��rخ8������1����"ԑ���}�Cc�,�V�2��� e�9��,�+��r��	�3��I�	�&�s���b;�'k��6��p�Ũ>0�O}ɶ��w؎�UF͎�;�C-�,��u��P�[�c�-,0 3�{.�������/1�X��+X�F��gvŽ>��f�u�O���O2�k݁Rm��܎�	u�����D̻HD���qW�a����~��䍾<������}U�������m}������m?j%q����������%�0f:9Sh���p@�ārQ�1v(/=.����J��H�p��C*��XW�vGu�D�BP]1�Dh�큑�o�Q�-9"Q�D_�l���J�`j�-msG^{l/��'��H�[?f#�������9��k�Z~᧎v��̨
at�Gn9X�	`�{Ot=gIv}zu�33j�t�'��ĚkLS|�3��h2�
"�pP��p]C�[c���P��bm�����9��:���M�9�������vu�$��#<-AP�9H���\-�J׽�	|�,DR=��3�"���D�jZ��e��I.��� ��#a�����N��;��aw	��hp�f�Y+wAYM����ؑqďo�B�ia���E$����0�haaٻeE|<(���@�6�V=69�_�zd*�_���j}ï�r�b4�a�W��a�3d�80��H�����'�2��W��m�JCT�|c�
x�g�kG�Nx�\���� A_\9��L7�v�&0��&u5���8����HSz�?��]+o�-��%'"Է$,̎��f�E�PHVJ��`l??8)%�4ƣ��k=��ԞC�%!�����z���4�tA(�����<�3�cQ
��?�?�&�@ףK<��qSVy��%=f?��,�0m�Q�<�<�5��A��E@*�(�z7�����4d���"t'��6��GS���3 $6��6��9�^$tMugw���h^zO;W�A�u�vr%�J}�m�B��<�{#�OV���`���&!r�n�I��E$��+�b
Vrp�{���J���o(Zb���]ӨV���ƄLj���__e�w�5b�-��)��r<Z����[�Y[Z6�_Whg;��eA����0�5^��М�<6���-/ئ'-n,�ʏ��la�aB p)��^#�+����=e���%P~��k������>�z����z�y�?f�DelJ�c��3S��ʷכs�{?��oGf���'�/���esymJb�O���Hj�y��Fu�� �^�&�Ih4_�§���4�_�L��Fs�B�U77�=B�#�֘�*H����!�R�k-e!K/�!�
$* �~v�\�ۢi�Y�-`UA���Hf
LE���g��~�ɬ\Κ����6�4q��]�+�2w��`0G�MN�	�eƲ�/t k5���Æ�`�rV1�2E��b��F�������)��H(��Z�mϢc>�ۆՄ�Pw1�T��Jk�$�-����>�ʝmk�v�/Ty��R�I�������/�R ��+����dv,�8����I��|C��*4����AsuvD\�9fo)/9_������
��,�Th�f7���׏5T��B��yڱ������c�5�ɘ���o�EQQJs�_�f��U��z	)���x�	YU�ok��^[��:|t�yS�N����GRx �t:[���N�Ś��`d�lr[m�q�P�+y�d��O�,��]���0��\2� &�o��|�#����n�A�����"~z��m^5q�o���&���lE�{c�g�z�c�-su�����<@�-�f������ z��)�˩t�c��� 6��ǩBc��*���D�$��p��I��R�����m�G��ID��!�X*y�WL�6�M&��Q�F��z�dx�#����ZϘ�:��i�]}s7�������j�3s6�G닌���y���Պ���dA�vH��yv��׮�� ��{�k*�r�E�)_����F�4���VRh�u���<�D4R����]s����k:k��.�|�$4�u�^�x��w�Sb]����g�1�$ ��^�A�5��,�=�Z�k8�XV���U6���%j�O��
:�˾^DW5�����,�7>pS!�o�dѧ�D]�z��G�6�M�}�LY9�b��Q_��~���w������� ��^�}���+ɏT>�D�>���|m)k1�6�N!$���q�#���f�MK��v;K2X�-���Ķ��A`�k���v��x���1�:��Y|0� ��Z�XH�Ѹ���VNA�aF��!����4fΤ�
��ɪ!^f�E�4Q�����O�F������2�\��+FXHLR�j@��u�vu� q!����Pef�]��>��i=�{�X�_Їe��$��{đ��C=��[�eN	���{�B�U���hH�%Z�n���%���Y�:u�9����,0�ʡ+�!dg �${��w�?�%��`�	�X9��76�1�\V�=�O�(���E<(�.�cV����ꝼ�g������ 7�k*��w�b��dC�K�1��[�T=H���g�̚���Y�Kq�
�Gua�U�l�xN�Ü�B�>3��_
T � �G���vkc6Ak-�cf�!����?��eP|^���EP���rMQ���*�o��S���G4|e�}B�)��'�+���'�R���W��������2���#��r?���뛔 L�2{.��
��	&>� ~�V?;L��M)��|�n�P���b��G�@��ltn�X����޻�(�b���uƦ�얿 @%Q�'9��n5X���%3�W�e$�X��f�6�+�2#�㵢S6��ߵEt��=l3����׿k�Ý=��C��j���U�2���IFh��y4�j�����,��+1nΨX{�<��B����?�Һ��
�J�LXlxV64EB    6c86    11b0��xَ���[��}P+SB���MB�Ąr�KY.��p��k��.y�j���C-]'�g�Ue�-�,�ZvV_~k�i7�C����N���2?�ߣ��AĮ�Q'��e�jW�>v\![��ݩ��"��[84v2�)ǅ}�9>taZO��0��Z9��?�e�?�7g�98=̫��4l[�ֆ$�k�E b��\&�g���*�\= +[I��yc��OV���hG$i���C����ߟ-��t�B��٬�;��⼼�<���<Oj���1:|y�,k���O��+�������t�8G��R� �+��88Q����ب�t�7)|<_���y�Քw�
3��Ҿ����	����$5=T	�t�
<=c�L�������*�cj�Xx �h;�<�O���>�ѭ���w�B��V�r��	��ԯnO���Vc ���ޡ��=c�\����V�r.?�)��;��]�)DB0�fǊ�v��S��g��A����@O�?Q=�Eq����?q�`n������T,��U�c�na��-�d(�/��C�@",���T�5�;� �v�$gB��5Ml��(^N����/�C�f9�l��.�r<�.���IW|:�UlI���\�x)���Dk���qǇ}vʃ�W�j8^e��8���Mp��p�"�C��F��.A�H�X��`�1��>���y
]������ޱ��u�z�dt?n�-��)uz°�z �P.^§�[��Z�A�t��w��@}]cd�j��r1K\�A���ZWm�7a�i�ډ��O�)n5�_��;W�γl��?H,[�QѦ;��+s�Lm(�c�t��y��0�p�N��Թ�i�{Dŭ'�H5A�{��ә���_��c���:��Tb`9Ko��=+ ��ͷ��y��IA�����'�Sy�R!F*�WY�'��l�:4�l�34Q���Y�B�G�Vm�B�'�&Z�B�)u{U{�ό�N�8��<8'�jӋ���g�$������˼Ae�i/�I$I1:4��l�����n8c�$�B����b����H��ͣ��
&tI�W�Ռ� C�H�[��LE��U����D�buJQ�\�#I�ײ8HD�v�\�z9���uǰ DR�J�v>�
U���"�x$v�*I��ׄ�t�P'�{y��6�����(X��(�<�+S {g�]&���D4�Y�9���͈�7�﷢U�x��������0�ߣ4r�@PM2�!��g8��|�7_s_���V�HG	�e����M[�JL׃4�oC�����$!7ߞki�K�Ɉ�Jf�ܤ�S,4�Դ+�����ϠB�UW��ؿ��=(���$�Q�7ȍ��3�ݶWI,��%�R��tw��yW[U�/�����(/`�e��8���T�~��D1v���:X������p�av�j+���u����ج$�H�-��D&/d|<���׺3��Q
��ɒ�Loi
�=yeЊ��;��c������ʸ��pz�5+#5�����,��6���������\r�Is����3'BR�"L�dNy��.���0>�	������"V?�A0U�;Q ����|h��V�(�u���64`��ޤ��S�B�j�O�����,cڗ頬.��\ӃO{,q���oZ��a��g�-����"X2�_�zP��&��� r"Y�	;��*��޼a����[l�SV���ΝsnfuZ�L
Q��X����Q�;�����mʱOx|�jhƞ`ւ�6֦s0�������~`�Kb�r�r�2d B���\�7�X2�։���5˃�-�Ȣ�U �bAZB���:l�^K���5��ga�	�o�k�U��,���B6��Y�C�]e``�A.ߠ�~��=�����ߤ1y�D�ZZ%O��q�Y%�#���,�4yqEp��"SV�"b�c�Akh���-��s��̋�|��T�Wo�>">bP�K{D�����
�T���+(+��u3 /�O�)���yxA�Ό!P�kN8̺�0)Δ�<��yL����^Ω���7p=?���eo9dĭ�l��dP*`�Y��'��X�f���*�2�4D��]SԬ�}Q�!5��s��-�y ���I-�)���R�>TJk���Q����T�^�JW�֧�v�E<��7����'W�BB�f�
'�eo!j�� )|]&%%��|�q9 I�;�e�`3�4��6���/�����t�	ۑ�M� ��L�=�k�=�5a$�#�(7�wD�RO'H�����I�&�EyCy�eU¤+�v9P����Ii�;�7��,���B�F���|/t�)�p�Y;Q�5�<��;"����i䤺������a�R�>R7NpsZ��{��{�y�v�Nu?X��� ���`��5��]�>N��`��]9�H�w�����S��;�;�~�W<-�;Q��W��)��aWh�h�5�4�M7���U`�1��3�� f�6��49�߿Q�T4ي�9\��ESx�fPtP'(%��t7������g��A���zb�w-������/��s.���'�/�u]�fUZ]{,�O���,��ء��İR�-r������{�>({+f�����Ǟ~
��O�B$��a�A��@����Xg��=�f���>��-*��sŭ�u�XGE[*+�uʈ|�M��ic�V��'�Td�2|����3�D�����[a��b��!�(Mw��Y�Y��ktjU^��m:
���FB��uM՘=��͟�v��G���¹l��9_q(t����D����S&�I���+��\�UnF�����.�P��n�Z�5"��ލ�iL�?�k����֖5�K��!:>��1�f�)1������\��8_ݬ˹w��� Y?S`�<C��3m'��S׳�VQ;��J��NS/P)�@a��Қ�^��o���ҡbOO2���Ӝ�^=�Vlҥd��7�"�d�8(�%��D��,�/��)�U֣�T�l��*EB�H���Ep�$+��`��+qHSC^���ʀ�����%�J��b��)�IGe��P�?C�Z�`�s�N����\��w�0��6��Jzf×�%1g�l��C4E��A��I7+ԍ�ŮEF]KA-
���,ѧW)�;y�.�<��{���p	-��b6Iut:��B�W��c����`�Ԉԗ.�UJ�:��F�b��j�����C`��i78�6u�S��\�R����_��*�(��	;6_��VQ*��=A5�1q�wA.~��}�/�T�D��d�NVR���T<��;������w�A�wa/�����O����SSvXlj��H���'\��$�iܦ�C�]�^����	�l7a��*����_��2%5�1ROV�T����e.L�;�5��"j���g�u�#�=������0�n-:e�98���I����IEw�}��=iu��c��S*e8��@ E������?�J=ɀ���l?5�����t�J�^o�a���WQf�构gv�5dT�r��7`b6)A_@2��Q�0��M5Q�u
��܌�ז-����Gn�R�R�������$ֵI<�`H7��k	���/��m��_�3����m�S�큥�]�U�vF�\���̨�cU�D�X�`��ߺ�1��%�P+s.j��e;��);GW�C&%js�a�sp�8z�.���1��N;��E���rzvگ����q��Q����<߳sp�]� ��I�d���7>GJ�$ؑ����� mػD(K&�w�~�~�+��F�8���(��V��g��L�A���2<l^�Zv~�T���<�ku��c��>�: ���s�RQ_�4�cЙ�ro�������L�� �^~��7�I�I�u������L������B���=�������7���t67.~�#��j���:�L����o0��0�Ԛ �X'8[Z_��T@����9ZbJj'��@��f9�r鎝�����{ow�Qzα�!?���*��p�çs
���E�7,^�T�����5�����ќ����� �tkNs�/)��zK�Jܰ�{��
|T�&��60�k�@O�e1h�H��Sθ�Zbm����=��s!đ�lG ��`�eҴ+�|���6T�h�(n�ҥ�5	gTH_�o���wu�f7���mRĉ :��O��Vx�K��p��Za�͗.�\C�0M=��u:U���{�˪��)`�,B�=h�v��r��8�F@����v��j�љ��?��E�;�y�^�&`Z	�|6�n�����'h$\Ʒ�^m
��7Zle��e����f�͗Zm�"$vH�	���qw�Ku@Q��X>�n�r?�<=�B��$�q���/w|ZxujӔ9�uE	j4�=�&±��jwQT&�Sv&ZN����)�r�����#]2){��[�'&\������T	)�^O�*+0��^"�eZĉ]xʢ^����Hγ���
@�: l]c��*jk�18��