XlxV64EB    4b67     f500f��l�j�K}�����sa���{sд�`�@�WYe�l��OQ[xY|�k�s��J"�C&�G^��A���p��a¨eƕut���@R%3����3�O~	�{��e%���Q9��%�)��%G,����(�װ ��>U3�Tv���A
�Sx��0_��Sb,�1��� �u�W���
�
�k�R��Zk �cu�w ƷѮ�˔X�� ��d�� z.Â��>>���� c/*�v�G>)��M#�V�m	"�N#�iM�Տ��T��Z��1qT�����Q8�D=�2}闺����e;vc�~Y�Yt~���� �$~����9j֔c^(�ѹ�x��ܞ��k�P�
�-)
NI��j�BL0�ԉcg���ͨg�����������3$�M:��u��a/�R3v�)��3�(`��n�$���+N$�2�E�s�ca��Mh����|�ŕ}��#�r��z:C��׃����4U���u�Sf��C}�H�|lD`�C�qr��c��0] 
S��>����P%*�}JJ��߷0����_I�ڃ|�K㑨Ҫ(0d�§K��NE������pd�����|��vo��tt54�a�5l�Q�A!7��+'�G��MM���9A*�	�0욳[���#j��L��K{^�OJrگ��F%�{+�2�\6�^`.jZV�v��ks�!�%ܭ ��(v�OL�d��"� UT�+]�w�O�^z�
��S��z� �7f;+�A�r�r��YG��߈���	Ѹ�Q.D�y2��Rہ.��z"��v��l�<����[�^�㎾	Z���O@G���x��1VR�lz�B���UY�T��D��V~W�o6�W�����5jAm��#ޱ���<��_��c v�";���9��:
 ;ݟ!�z�
��79?1�|�HU6��uv�ˢ���Lc���f��Y��M�}T����.R4m/s"�©�����ݲ������KE�퉕S=M�~G�R(gM��!p��-y�Qy�QJ�
�	u>�� 5�K���5~[�H�����*���0����������͒�_h������W�U�eҜ���Fn�S&q}z�����T���r�j�2����`�P;��xe�!i&�1��qm�8M�A�u��@�?5�iA���߁[q�������3 ��� B*mFݱ�Ʀf��Q;�--8�Xnr������Rg��Z 0'��F��i�-�Lw�J~@�m(]�1�U��>q!�*\Յ���PvQ��&��W��dښ1	�,\U��c�s�&�X�L�HF��i͉W?�KH��۔5<K%�q,��X$��׋2B��=��갂��m�}����u�:һ�n�{^�s���\Y��~�p�'�9����\M�6�
(T���~P�nT�!#�Td׿<�$x�{��ԁ�%j퓼��rS��}�[z_^��@��rO����#��V����D�@:Te@�B�:e}Ū�䜏��U���k���ɹ2e��|���E���ƛh6F��k�l���D��`-S�D*�/����c=s�M�h}�Hr�~���b���7l;�)!y� H$ܩ�K�����g�����":���</5�p��+�6��~�JG@���D!����.9�8�\t��(D�e� 9�Uua���uZ�ƅ�sEm.m
�_t�i�[6��D�۔4���f��X���)�`��I�`Qv����5�ꝸr13�|�eQ���5E2�˚��(*�v��D��|�En�U�^�Fa.g�ĺ��4��Ӯ?�2-��y��)�Ë8��i>WP��a?���]�|�����W���cJ��*���|���>�fs���c�������T���J^=��ڄ0XFו�/��M� �Cͩ��a֐D�;)�)�^��hO\��[uo�z~��̢����J���)Ɗ�Śݺa<��	0�pG�#����8d�bϜ S���D��஫$pso���MF�@�~����qW.���x�V��Ĥ�p.��ϭ��/����0X�ܾ�hC�b�SP��1���l%�ǲ�w)�	`�v;��m'�$(���"���L�|Ҫ>�J��f�q�!�a}`6��(��-恱X�U�����o�ӗ���S�$�Ȼ����w�Ϥ�U�4�m,F���B4��q=n��,a���.����d�C���2��`�I*����˶��o��cV�$���2�_Tܶ`��ig�Ke�'���c�*��,'��.�TF5�ǭ��+�Q~��Oߚ���v�G�Rc'�6�����3!Bp�!9_�֢/z�Q��u�Y��8c�LL�\�L@���pcO�4�������,��t�v�0���o��(��,�2�H�m7����և��K��$�p�@���I-s�M@�:�y��?�t��6ۡƞ����g�y'�m3�CQ?hJ���F���vw_��O�(����۬
V�t�t[�����?��zѽ��1��(��{#~���<s���+v؋��Ŏ���qm�%�[׈d�{�᫞��t��"��D�)�{��IƟ��x�E�p��<_�r��>�-o7���7�����z���|:���K���� 8�{��Y� ��l��.���g�[��^�Uٞj���@4�&#Y�x��s�����R��-�iw������h}8K��VF p�'űgƬhCq�	��3��rW��������������0�5�.�sa�rܖ���Fb�l���Q��E��W��sm=��P)G�&�#i�Tpw#�U�^�KDe$\ȀTM�m�����ߦ2�آY���wAi~pdVAAYy��γ¢���\�;)��J���,�9B�ӣ��M7	<?���ڭ�x`�z�P���ѽ�2䏀N.wp0�(sߡD��J��;���S�2��>ϋqe5O������.㲰�x������\dkXj�v��2beWk偓�a�vq��( Ѣ���s���q��-���y�Is�ض�����M����ҋ��w��!�C8X�0I�OG�Z�scG��A@Ru\c�	'�/?��v����1^θ��j;�# ԯ&P��(9���\7�k��"kiY��,��D	��<,��(>t���e��C�9ՂS.���X��#�(�"{���Dos�b������c��d��J�xP���4���������x���E6@��ת �c6�ܗX�kh8�3W\l��C���	َ�'_j��pqdq��1��Ax��R�q1���bE���4�<���2�i�� �ܻ�Z�[�%��~�+;z=�'�[7����7�N(z>�����L�"�h��
��s/����EfR���:���kL0/(�^�P��\N�!Z	'���3F��X�}p�+�m�hT�))j���(L8M6Bz5�� ���g§� ���HagͶ���j�Ɲ����V�e�2��cʻ�0��D/.�q=��Ŵ��xl+����y'3�L�z�&k���G5)�ID��U��S���+�)�)�ލ�3�%ծ���Y��p{��+7��1 ���+,h����r��Y�����2(�_%�@5��(,�!:C�11?r�#��BU��Ow�gz�S6a��kn|�!�����)����/} {#6Cڦ�W�,�%�~�,�v�#F��d���zG��j�A�'3j�B������Ef#��8B�O�30���{�c�U��:_V}_��nL41A��]��KM1ۥ��W�����k��^Q��)xo��T s�@O��_mf���b�n���L> i�V��{����㬖9 >�ێT@��ri��(v�4B�'���Dj-�+!���