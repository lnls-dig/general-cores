XlxV64EB    1ccf     9b0��=\�TX�D
_5r'Uvs4�X��yXyx�)XU��b��,�;�5��&��O�T��a�m�8Tݞ
��W �	%���J/�)�N�`�6��H���1��ʚ�I7+ƅ��c�~��eM/�UWS���+1��,e��l@ ���z�4a�]׾c�X��(�`�V�T�����gH���r�:L0�֖}Y�"��*�0�h��i��^̌�6���z]sM	��"�D�)�������sӛ7���p���p�3^��D�tι�e�r7�_*��!�4|�1���C��5g��N
)�(^��kj ����0�y5ceaP���VF�z��7����[�A^�����|Ӯ'�h� ��M󇒧w��Щ�������k��Q�0I|-�BoA���ۮ#�񦫲˨n�׎̆ٽ��z~h6av�x�>䂥�V�����d�a@�j���
ib�K�`�� ��n�5%�nTs���CL<��FK��q�<a*h�(�z3��	�k��,!s#��>c�c�G��~]���!���p�x�ۄ�O,V�N�7i	8"�DY��I'\��՘=D���Cz��DsYH����`�z��h[2��O�?x`Φ!�sH_�І�1�,@G��9t���w�)��%�=e�ŷ�A�8'��ɋt�[DI���u�A!Q����o*:����&SM7����S�-�A�tdkΧd85�[�xg��&'kL���ZF+N�]��Q�q���JA6�ϜW^+s���ה����"H}F��y5�,�!N��F�t��{�H#�	��s����rO��%�ѰǇs�}�A˖.{S�H2��Vn�V���)�5B7[p�t���*�J!v��LP:��v���@ �}c���ni�N�{�c���pӘ_l���<�֨��_�����/�g�@ɡb���.�-+#er���Â��B�ξc֘�o����:��|V,�>N�L~��쯫����፤ԭ�2���Wg����x�b����(+ʾ�5�-��T\��`�=���׆����ۏ��<)�\^�ƂQ��vy%���`'�邍a~��]����*/�
�Q�e���/K��I��I��s����p�\���HO�X�����ۢC�H�sE��~��-��ȹK��T&���Y���\�b��1&�	f`��"�a�>�C��&A�!��vJ�7p\�n`e���(ԡ��
�]�)'H��|���Wy��򥱑c�l���L��h�ڂ�����{���8��B�E�чF����{�����닽����
a"�R�0��TOE��"��1���U�I]="��HP$�f�9�O��''�_t��.�7=YD4�k��>�F���.8YP�/O"�`ޒ����	7A ��|l��*>�$en_���q��;�DX�每��ȼ�O�Wv�h��Q
��?Z��~9i�Y�8
�0\/�V{�>w��[n�w�w�槟��cE�0K����_1�ѝΊ�����XȞe���b,���j�\�F�
�!�4����Β}�7Nn8��G�FϘ�@ˋ{�G����X ��1�ߏ�"�:��r*��ZdRW��o�0���,��j<ӿ��2M��)��&bu�ꍎ^�}{e;�>� �|BN�[�⺄wX��/���Q�`U��Kd�\t/5�o�NF�j��[(>M����weYr]_sC��nZ�&x��ӌY���D��i�>x�ݤ�s
����J��a�����D!c���BB�P�sh1�p�������(B�	�B8x�d;P���v*�fK��s^��e�H�fS��TC03���q�A�F�Iβ��K�l6W��͚���Q)�O��@�5܈Lmzb^����͆��M""�,*�Q3ӽR-�g���9��x-�v�:����p�|��\ơ���HgI?7t$��2_��z�(ǌ��Gk)�G�;R�]a����{`�!�>p�z�ДR�~(��S��@3�9��u��BhK�$��S��kk�V�xy�Ho[�ج�e�ϳ`3�J.!��%r+��L-���@�|�dsp�d�����:z���E�d�0����k�g��������v�s9I����_��Lt
�b��p���傇����W�&�G�=�Tp?Z��SRIv������k:a��O*G��n��_�)���)��j�&�|l�R���w(t#·�~9J�ݓ�@��W�9�	P)��BB�Ѝ��@��I`:���GAAGΨ���X�êT�IL|�����|��K$�e�?
$�"c
b],ñ��ل�(&�/����>����'f�۫��VW�A�l���v�B�ڭA ���h ��/��Ԣ�t���!�/��^!�����ǫwR˖󁵓��t����TdY{p��&v�;U՛6��rp1w5t�g�4i�AL��l��cc��k���0�� ����=aS��~#]���3����2����