XlxV64EB    6024    14a0"��P@[�k�����������j��v�C����۔�!U��P�ɬ�jٯ!�ef�ý��m� ĔM���΄I����oh���խtW���2y�,���x�fi�o�+^H���g��$B���(ۙ�n�I�@(�E�К}���e��=������w��Rh��].��Rs"��"�f��a������=�^��?!�(̋V�,m���Y�᳕��(o7O�q�d�S��K|���|Ԙ�)6^���Eߥs��n-
�L��!f��Q%P�m��;�Q����G9�[��q�����ٕ� �D��:���-H	a2�>+�/TK��:��`|�E��T}�q�U��,t)�_��i� �
yH�/��O8��w�k�����6- ^�������E�.�-Ŵ�¥|wxԀ�a��t����C�{_��4i�E�����Ӈ\�7�b��;�����b���
��O��Z�Uj�X;���cIK��}%ږ�c��
DFM���n��Ijc��Nߴ��JE ���3 C��!�Kh1���b�u���h��9���� ��H��^��o-s��F� ���#u�)%�E"\�b��<��k�v&^��9=�\w�0�X�������E&�Uf$}��x`%�y�`�o�eW�=ܢ�i"��7Y}��-�Ӌ�(�Q�#��gb��Kďm�eWB�����1o���+�P���盞�˷|������SM�E} ��K;�N�}�6�����\ܺ��.Gk�8� U�&�]tΝAﱧݣ��x���;ZW\��/�Բ�Ʀ3��ƈ4����Џ�š��G��ރ�ъs����r���[,����6Md�?>Du"�+���d�D�׉� X���](V2�j���x}�"[�CD�C�yl�dT����=��8n+Υ)��)H�ķ������u��9>����Q+��X��t[f�Z5]C���O��雽��4��b�ȅwe��k�z*(��Q����_|����b�����?�%�\9�^P��lvGڛ1}�L�i�C�8��[��$x�����~?��'���4��<{���/hC1��� D���m���ė���!�t�t�q���W�>~RS�c�e�a�?���4��rJ�~�!0�A/��ל��r���j�5�!���X�H�=Bi�!kQ��m�d{$զ��i�e�!��^���8�E�5��0ǜI�d��Lؐ{�T[:�H��٫nT)ޫ���6Vn�6zvw���ݕF�pԘcG�0.�+��$,4\/̅~��"���\�IW��� k��.��o��w���]�1/^����
6gJ��2�|��_1]>h%�YK�����#�4aӁ�uu�C�p���P){E�q�t����զ�Y-�3�����=a�Ճ� A�`���ءJ�� "�3�Dt�	�dg/R�(������[�Z
u�D�N��ᦙ�ot�>D�Nx�]8D˳����M�V�9f6	O�p����c�⚩��mB��y#�z��������g��L��ĪsՕM1����	tRR��s��k5G�[��!4%R�C����W�S�Ʈ�ӷ��v������
�:l�(P�e:B�I�U�$Z�~�C��R	F���}��h��]_)vZ�����1w����K�2䊘�@ߢ�.��ȃ���\�F��)�a�݁��ll�.�J�Zr�ndI9�X��4d�#N�.��T�F!��bI�P�g%�
���3=�ü��DW�/CZ�.�q�P�ѫt��jw�v��T)ɓ�7~�����W	�thym��P��3-_n�Q��aᘓ�Pz�����`ﳘCeV���!�)�W
aL������9��N�l��,��Q�C�uL��Z��_FRZ��5���D���NS��
v�@��s'�+q� �wV%`�Z��@�	w9�UK�T�~9�~~�N���cҧdN:D7 V��w�7
����_ ���˷��4�i�`��Wd���ԅ;3���v�Z������PZذ΢�$k���/m����Ͼ�&j��JV��϶t��B2).& z��	{(������R��Z; İ�~��]W�~=]X��4[PF������q�W���a�Lh�Cß~F�Sx��|�����4~�;��Z<�_P#�'�yQ?���>x#��=�l���cΩ�C����G.Cm<�85����m]�mJ�|^�G�R�ɡ��KHi�xtƘ[u��v����
���f����
`]c���b4U4�
������ �����UT���$�e<��lV�Y��"mSD0��K#כ����d4���kBnhIdS��m(���y%����îG�ℵ,����d�*�[lE���X�!��F0÷s�3a��x��Lbs���m,���lV��J�5��oOfpt�2G*�k���y����Q|��1���$ᣟ�ƯƧ�̗=ݜ>������:��ف4�?��nI��������������ש^�}�ӿ
��^(�H��v n�������Īݧ��[JPzMux��t��m���E���E	��T�X}�9��ޗ�=�uVD�{;j�����v���& ����ǯ�PB��nv����f��J���d�L-�Vӄ�J�s�[�
��w3bQ
Y�:_6]V!��f]�+�Н�p.v�k�;A�2�%V��fP���o��ܤA���=r�P���"������Ǜ�aj�
El��bLբ��('P4UJ��Ӑlb��eYd��h�F�?�0����h��!�"�B�4��>v_�TՇ�O���)FR��&��e�~_����.��ZT����b��+���p�Y�I�7�uQo�8���_��@�Ż��.S��th:ݞQN�)��^�b�/AmAf&�f�l��������M�P�JL(S��U3�jo����
x��ݼ�D�އ�#���oI#94+�khsz�����{ȼ
�Bʖ:�@a:����M})�Nb�ѭ�D ����M��~�g�)����t��9��s��}-�͔	�m�9m���@�C_s>��g"�Xi��X*L��,AXkn�����K��^�aH�����}j����m�z}٢V��,T�I U1JTZ����I%���Ť���X}r^�?�#�����x�$�,��aAA��jQ���Iw���� �չ��ϼ�e7x�;��Vn�4T�pR� 5�}"J�{!{?��6,��P��a�7(�N��v���]}Q�������o�~�F-C��l960M��Oo�Kٛ/c+�v�{8s7'&ʇ�B�o��p�C����Q ���ɕ�Md0@#��2�K�S�^��}ԓ0�Q#��C'�ǫYe��P�yVw%�_t������i-�^n��<��,Ɇ�+��}:��Ѥ��� 	i�jZ�O�	3�[X�E�*l��8L�����^yR�d��w-��u���%I;�0W�2W�Dʱ@�����Y�����	����0(ju�t�o�kdZ���R��ouO��:z�k?s�fl6���m�-Eō���L��s��sӳ���Q�{�L]6�$�w"�!���D���X�ԇ�X�l�Ѥ	v;����~�[�Z�8��Y��Q;�J���q9�x��p��M	cu՚�68��寧?���U�W�I�{��\/���-0��b�=��'�����"��S�Z�������	��j���?n���_U���NL3�X��=T��y��;��HF����<���[��,c.?9�E�8�(Ae!�T��d�/�xS�&O��	~���g���DL���y)-�Jq����P]*��n�s�EL+=��{�D碙��Ac���j�dEDm��k����������Z�v�<�A?S�������4K_��jT�\r}/�M��M�u\jy��n����*.�'�����ō��4�Ʉ�:����.K{Pl!^5B�u��>��h�0p�<�F�~&!�<�C�{�r9��a��!f��a��$e��F���(v�D΋��m6%�K`ɜ3�qS��+�����^�.�(�@O?#�щsc�����/�����-��[����K��2������!#ﱳ�csT�,l�TW��01�>�E.s����r�I1mG�4���<�PR�c�H���7�DvzO1g������u����B��	_�a&^�q%`<����s���xX~Qӛy�e(O���"����hd�Z�~M�ge;�(F� ��5�|�x޹�[����΍���%��e����rɽd�Le`�D��gU��<�a��Y)�{!��I��h)����y8���P>���m��\����aӄwz&���5�/g��{��z�s	< S�_~�~s�:�C�&
�x��g=@��
'e��k�9��!JD����ę3�4�`1���:~VL�vPj|��ĵ:a�ةO�M�e;^�G(SJ�0�@�A�b8�p�9/�v�Zm�!ɾpJ�h!���ӃԠ�~;I�s9�㤠��A�&�ZGM�{g��}�=Y(���\�R�.y�n[z6z�ڙ���؈w�2����%A��%�I��I� Ɗׯ�D����4t���-kZ�����8�j�ȣ"c��Br^ՏM�a>�b�����,u濚� [�Ϻk�,��l�`c&:2�k�Qr���O�iB�$�t����Byr����@��N���^e��r3V��Z��������I^;H)+�^�L_Rr��b*S��O�~���	(�>,Su�yosb�����5A�莕?�z3���4�����ĐHHA���:�i@5�u1����fňڗB�5+]��i�����!T�`��X�_�{��A�����Hc �������Sg��,�1�;s�ٖ��o�Q�kk������y��� ���'�P��L�Rjt�2���5��S�h�֘i�>^٥��y�7�>������Tk
s��K��ox�0w�L��|U�_��M3yD��;�9��/�E���
�$t�v�FܬW��%���c����6�g�G�W�~n�
4���Wcp]�z���+M�$}e�٦�����k�\���C���	,�����4̝�@���?n�cR�o����P�c������ѿ`&��+
2�[.�� X�C��У�.�5aa��<�v�������3 "�˔-��B�yz�Dƶ��
z��T�F��z�k���OY3=S�VI�ρ��>�5��b��B�P�����/