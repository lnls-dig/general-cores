XlxV64EB    222d     a20�n݂�to�X)���l��O� �s�F��������l 7�q����ˬ���:ʘ�9$M��J@��R��p�|�4��Q��A��:���������?��a5̱�"m8���牲l�Ғdڦ����œT��`� �i
���9V�~�4��]������K~���g����^3g�]�/�W5��;)	
}�t����L�Z��x�d>��s7�2<��O�<��a�3É,�|$A��e�W�F>}2؍����� �T�i��t��}=��� ����w�l_,� �[L��6�+���ߟ�~���_L��4Ǖ���A,�&-]�ҏ�W���ɧ.q�x����K��Q�'��Ki#S���#�4�`������L�n�F���fXn��W��)��+eLH���2M9�-�	�,�JrO���H�Y|DH0@����#��6�C�.�Q�d��D��-:3
�D���R3�^�����;ܪ���3K��0U��8�"�a�9��TD�?C�l
m�R!���S��u�:'0@�Tn�M�(ɷ�=�!����u�Ot�wi%l�i�cҳT���#���ͨI�!Ar>DmTe���<�qv�!	� �zI��<$�|�6�y���4�mJ!D��D|�f���w���
	6�-l��z\�/lqӮ��YȴK\)��
��4�$K��,\"/��3��12*�9�V�M��_&+���Z.j����ʜ�\��-������� G�;�9�Y	��'~�4#k4m�_��:
F<��Z-Ȝ5o�X)�=�2�����E��i���X�
d���;�C�3(ߪ�b�����w��Z�)�W�¡���5&\�!#�p�I���fHy��"T�Z�<V%��\�����un��FK?L��s$X\�z����P��'��ucc���
�'���ұs��Z!�7vq��Ufռt�%������Q?�v�����WǤM��T�)/�^Y�ߨfo�SN�/�ϟ�k�?�va�'�����l�A�$2(`UBк��T9��9�?�ϝD��Z���o;�J#��p�z�����Hpy�W�'�O��H�={I�r�!E,Wfpsd�����}D�O��B�V�F��������=^�"G��v�~�M�ᚰp������#8��H֗�C���{�M��a.�|2����)��l/�I�4>�u�*,H�F�s�T���\c�H��=w5]�3n�AH�䣁���/�l�$'�E3�Փ9|c���qq?le��"3)��_ҙL��"���
#���G>��fd�����D!�v_�E|���Y2X8��h����\ʵm���h,L���fH ��%E ��`�v���h-} �T�"i��[��j���Œ�ϸ���@�þ��� %T��i�c�<X+�Z�n��(�D�v: �����(ayߵ�����T1:��&g�Y^����2�U�L1������O���ۡ�>�,�~+�w&�At:�D*�z�(���4Mb��v�vd2G(��&&��DJ����!�r�Ҫ�!�Ga���s���+J�������"��V9��mu����{9z�ķJ�qL{ \�#���O3��v}d̌��Eo7�����X�|B�H��"�1(J��5Jno����mz��l�_�f`G;7VQQ���B.5q4�U�����ҳ��ccs�1mv�{�_��Ĥ���u��T)?�}�:�G�`���*;�7�/� g��J�W�A����Li�;9�4�%����r�+���E�*\��e��]p|�
�>��1*�1`¶�m6�����`�'�E�ju�sו\(6�0��pڕ�A��m�� Hǎ������A6xaT�8�.�a�CO/�3á~*6�ө-7�8�~<&-���EUE�
:�g��λ
�og:��Zì����-I�*��`ً�^v�
?!�5�n���A�Ҭ��Z V��ݼ�Ai\�e%�.���F�k̦[C���E���C��vk�ƿޭ�C����k���E�d}�GUDQ�/TKĨr�t�?t��Q15,����-_����jG<r��$*mق��G{	~�Z<�Hgi��
��ݱ'0rX�0�)\�#�(16���^�7ZH%D1���gW�P�.�z/�qS�uM��$R�h���8B쐯8>`�_�{LO�3��5A&g��M��i<�-�$���+���*O���W	���z ;�����x�H#�xa�����T�m�.�U�y`��o�C~C�d��XN����R6�nζ{�j�d+Tt�LX
F�� QX�E�ml�P��%R�!õ5�S�nl1�����*���N�2E"�=�i}?��(i1@`a���'e������寎1Ѽ��4��N��:�<�M���JlJ���6`SH��v��ˉ�6�HF�&���a��UQ����{� ��z$k0�(n�uЙB�^���A�S��y.
Ɵ��JCL��\ε��?��\���C 2���!0_���Fh�8�+�O��#I���rv_:b�Y�S����K��X�~��j