XlxV64EB    19ea     890V衙ǽw�fY�=Ot<`u�������1/�#5�3�[�։;�)y3��t�-3���.�~�Тx��+^����7F��N�p��7�Y ���x�=_����=bs �`�|c1�� ,�3	%�_�
��[��GMu�Wy��ժ!:�j�`���ִ�2�/�wa�5��\q��N��o��eeպ��
 N�g�tݻ�ogM7J7�T�.���ӵ��"l�����=��}Ɣ�3����y�ӂ�����MȺ��ҳ}��
�|,�p�b{�׼?��'5�R��"y�'��~��[�uw(;+��rxRƨ�2��c�/#�� ���x��}�{/�yt��=�}Oa�G]�������ʠt�rgom�.�H��K"�bł�Q���^�)@�k�Lĩ����P!�+^]�m9՝&��:�p������8���W?�U����J��4����RG��-�븷f!�=��N|����8��FL`�u�l!މ��͎c�����F^�P{�%�����&g���H̿��;���;1�a�M�~����]���%�Csd��e,�N��YyA��N�~��lI��W.,�6TT|u���.�@D���wu��q���H�}���?7%b���ܡ���zr9W�4�"ZZw)� 2�֌����!�j��D�v8�%�ر�B��@t��z�+ �ix�YL%Eؖ�ه�-�a�4��Y���?��r,� EC<�µ@�3�z�1���%�I?{�S����=o�"yI$]7WPL � c��}���~��wb*Hh��1�d�l�>�z��9�����7�x
�D=���h���F!�\�ʣ�jvξ�k(�En�=	�qͥM�-�b�,��6��zC-�U�?�0�k��=Qg&�C㽤��n�-I�:*�Y�h�!^
T#B!���X���0]?�3��iSu��V�][ݙ��I�+�J�V7��$y0"xP��I�9��T�s�g��b����eB��5��]X��쫦؎:?�F�ά��*���EW��1)����Yq��cg>*:�@T<�Y�#8oJ�1L֏y��*�;ށM8Z���u$����'�ӕ�_�5�=JJ�4������.T����&�/?���%�p�C�	]|'©��$>�P����~�|������h�vP��ؤ"������6�&N�\�pa>�}����:#�n�UKXb���,�?��b;v8��ț�g���L��Z�2��u��uv�4�J�/�-�
��1:o���{�U'O�>���ޭj�:���I��;�Lg|��� ���հ�}�e`(HlC����7�qN�e��?����}�.1:a~���1��l}X��x�5�,6	�!�OZ��~�eqW�����E]�h�:�0����Rr�W[��`�?�e��L��A~�>��J�� 顚�t����_���Z�l��HjV��T"��7���x����q��)��<�S��ɉ����]	�u�Y0AS��!�u�-W��d�q�t��	�v V�l����Ѣ0us�3n�D�d+!TՄxzR�����~�S�r]Y��#F�s��f_����+n�tn�!_Ů[�7� �\0�8��x�Y�3�>�o$�2�߸�e��$f,۷�7�,�KT"V�;��-v��7��Q]��ͺ�0*yd7ZHN@��%���?��+0>�Z�XcIX���Ǖ���psO8��1��^歒}�ٯ�j	Q�%�.�h�R�E~�HO�n�Zxf��4��O��������u�G��� �P:�>��#����PC�.0�;���E*<G��z�y9� ,N�C�+M�?A��������L9j2��Pl���p����8X���/?va�>���2f���d�O��������M@����wA���n@�v�"\��!���u������.oh̊�BP�O��s�lF���Ʉ�v��>B�0e�`��2��3|����Z\-b��[����z�++����d{�<;~�U�m�ը��{�b�llm�mpQ���dGp���Q�������|̓|��w@�[*L�*�	�/Z�Ɨ��7�"/� ӳ@��3�f����Wܹ>��(N�o��-�����t���o�ѦS�C��*ԥNMZ&���!��u�f�,��h�-�?���'���)�N�>��