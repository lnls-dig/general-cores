XlxV64EB    5254    1240���Q���۬����PR����yl�s�� �Ds2p���$�2ϻ���Γ�A���#�� i���l{SM�<�$k��bhp����$�>��
�QÔ�����}0ruy!~�!�5���g�$k$6/��r�X���a.<��lRk`������u�3�)�tx$r�Ы�d@6��f�V7#tA�'P_E����8�t���*;M��?�Dדuȧ4�K��c�MP�er2peA�K��7���rFCu���Sb�
���*h����Kn�έ���/��� ~��j���	��@f�ɸ d�lu��Q�ǘV��%��SP�1V�Jտ� �U��s�XM�/��ۓ�گӊ�H��$:��������>0"`*O�o�ZAa }0{����
��_��z����$�\��7
���\`����f��Y�:}�1p1���k���4���c�5��r�?���z��\�Z#=W[��	�V\@)~xx�#a�޹
g+�Js�nl3�	A ���H!��qq�#�vJՃ-g����T��_"bg��M3VS+�vy��m�,�~T��[��n�c�Vr6}�@d��� W�+7lXfL����6��� ��`�_.�ZΒv�]����ވ��a�����Aԫ�^��������J�F�# uUe7S��P�yX.��Ʊ�GO"0�@�֪hԊ'����"��[7t��Zf��U �$p1 !��ś>5t���G�JQEt&�:?��ty{Y���_�V�s�{�!ۭK�d@�a�.�$X.L���_MO!����<A0::��`)1+�� ��A?�?��2��o�6O�n�G�#׆��Þ�%%0�	@#��[8�d"[� {��e���kjP��������\b��kޖ\�S�=Y�����d���_<�ȥ��"���N�`��	4��pC���9��kЭ,�fMb8NÐm�c����?H����_�}�-X������u.З&�#4$�X�1�Yy�vݬږ��0��<]$�j4k[���8'v�����B4���A���i]��50��8�B����1�ˬ���e��O!y���]�r|��Ҷ�;��}�F?�C�����T=�~�
���^�ʈ�rG[� �u�v�=�{n&q\g7#Z�������;�1���hK�чH�\fx��c�?��Ί0�D�G%2^$�e��!mx���XvU^����&l	�:C��'����r5��� W�lv���g���9W����NL�:� �9�ݮF�v馄G�7+Wn:LM�p�S��]�&եsQ}�U�b���SV�+~R�}�S�ͮ~ X�k<���<1���-鿁��i��� � w��+�.]F�)�pb��`)���~����i����rzM����&��2�=;�:�چS�'���O�G��\D����[�����KjZ�;�$V���ڛ~N&\�`ݿ˄w>���)ӝ �	�2n��Kڥ4NӀB�
�[��	:�F��K*8�_	���%�~d(�[��
Ж�@p�.� ��j��K���Ѕ���6LՌ�-���&C�#I�7Ďù׬�zNGKRٲ��'��>�	j���^�:t�N��Lsm���b��6i��m[vAN��n�l�$xB(��N�A���ǅ���֑x�N��{�u�O��S��[H_.�����1:�oW�a���U���{�"�u�c�&@F�����ך�W%HI_��o�8���zL������髥X��'�v�`_a"e\
X�E�;���3Qܴ���+'��a����DАù<%8���ȯ��+9~)�4̒�G�Ĭ�Q�-k %����[�-���Fq+�flA3�>��%\�"�f�ɉp�ȶ���;� �ܝ~9*��o`Ys7I%���!����|�OI��U���'�$�V �Q��������?�ɑSY��W�����~"��jF;(3��m���uZ�/�U��z��c���Y��d�f4{��*�y�R������e�]E��������r�=V��BTW��,c�u��3g]�I�BDW�QǮ(�9Ý�qbBܮ�"��rĸ"�W��~�^�����=�`ŖM�O9���sa�eS���K����|.{��r��խ���
�"n�W���i3����yx<Ԣ�ΤW�:Z5���'$�&у%�MPr����Z	��Mh8�W,}�����n���s��"�l�P���֑����,"X��.]"�A7� ���X$�e�XxDlh�`Ix'��&N���EK��so�t3u_�>��	$�ۧ���;r���=���A#*R$�ܐ���DꢠY�Հo������u��-���8Gs+��"�љ��Έ$�7� 
`��N�e��ӘK۷�8Q��c��xr0����h���+Ǒ鷌s�i��zJzv�taÿ_k/.0�m[/J�=�B;���8����qZ1�XcqU`@����J�Yw���� ��\�{ k��;�"
&��`�2�V(����b� n�1(S0�nt]��M��l���(�m
j���l�V��p�炶�
S�*���`=�*� ����N:�3�$�y\��~[��KҔR[���K��&�7���Xrg�/���>_d;&C?A�=�qr΃׆=�͏�|��w�ຈQ����̆if�]e=86���4@;1w��ה^�����9���8�s����WMFaVV;����]@^Q����FXY��6P*��u��YiHZ�Ѿ�▙���]z�TR���ө�Tx��&h�bMY�u�����p�'6�.�I���õ-�d�~MI�_66u����ZH߱���~�w��D;^H�{���F�ϋq"��3ۧ`�B[� P�U��pۇ3�4�ip���86�Vw�4��NT���P#a�wOew�����)+�s�-T��.�Ab�`u�1��O��s�ʨ�C~r�6F��q}G]hr��m���5�Myp�__�x�\8���ʜ�~�"ږ8��?h��5y�xb���I�ZbO�Ѻ;4W�A^����+���� ƻ�.o�����>>xV>��=_ntG��T}>U5~YD u�q�������Ea�$7j��)�_�x�7�7�X2@p�>���%Tj��)f.� �5',3�ù!��JB
�Y�iz�X��@����GE��"���U[����Apoj�']��q�����{J$��z�;4m���1�7�9��攰�.n]�h#�*���i��#�)$� vlH���M(�P�C�&�CW�Ƹ�v�.X6lQ���#؝{G�[�I�2��?:��t����H����B�[�R�H?zosV(���qۚ�	 �O�~��1Jr/ef^��V�q�S���f�F�{�l< �DF��V�Kj	������J��?��~<4i�����|_O�I6u2&��k07	! 7?��J��r�xI�?ujH
��|���%X��c���+������u7��@iʫ�k��E}�����9����\��H�L�ӭ�U����v�`1n�U�q<K�g��Hip̳�-Pu$k��l��0�wjVݘ�M�%A�uX/b�Ƞtu�"{�B��]�C����C��z�����/=�{N(�:���Ů�`��?��ia�lL�?ی�'S3��Ǧ>��c�n��a�rf��fbc�h��S���L�8�}����h:#{��PRE;-��m��4��͠"o�0�b'|��Ѵ��-M���ᵶkg��9NםSs�>3.���r����2V�ol��-����	�����s�I�c�sY+9RO�)��"$�`��>�E�Yi�]��19̉�!�޼��o�K�q�������#�IH���:�n>ʈ*�����S�?ΐœc1�@�'�''~d�n�L�Q�H�6��T����h�D�mF���f�9e7�tU�l_�#����ֱ�c�N�����Y#�k�8�Fh4h�7 �G��Y��^s���`QI���ɹ������?v%��g�>�M#��;%_C���/q�g����*����"�Hm�#*���!l F��3��`\]��{[�^��rr�v�T����/">s�������~��
�mC�Q5�q���5�#m0{M�Rk�Q�T�]�����W�Y�p��J���HF�N~f�;n�ޏ_W/�n���!��^���+�.��A]o��Ec�jM%L)�$ڬ�8���+�3�zBd�)-�{6j]:徆�/��'U�ԋ`{�cZQ��ml���IG7hY��h�-�/�9�'v �,�<����N����rO����DBj��>�ΈO�T�)#�U�z�pa���~�P.��I7ǿ�N�� d�M�0��+�3��a�%�;��r� �����1%a������g	���qk޴�[��W�h�ѦDeH��%�����}�����.D}/��}d�����r(�AZ������_ܴEu�����O[Z��v���<�R�?H��;O|X	���'Dhl��E-@A����.2�FWZ�H����yÒ���IT=�����
ۆX��>Ɂ��%�cߩ��[	ך���o���;����N橯ffl�L]�-H����~/�\ƅ����	��~˻�