XlxV64EB    fa00    1fd0��ZQ���lf��i&{���\���;m�)űr}�Z��@0�T��Nc��毷�߄��x���Ҟ0B5W(�>�w�Ȭ;ؚkc�{ܴNP�����jC)$��3�&��A����h�d��{�V�(���F�H}�RN�p�vOm��AJ�ҋ���c1��>e��3�x܁���V�Q�(-�2v�y��ӥ&

�%�� (39�E��l�[u*���R��q�Sa^��r��w�H�5��UuC@�T@t��pm�h��u
�f��]N�g��)�m�ΐ}	�.�.�d�F0����;"�ȝ����G�E�"�7"�:@FE��:�	�����CEٖe�d��#_5��<���T@�(dZ��&����7�ת��X�䗂Jl�W�A�O���B�[DO,)	x7���aQg��h)cV�Fͦלm��1C����2�d�\a_�n6k�;�8b�[�@YJAY;}b~������d�j-����;"�z,���'�
���}^���=N��.h�-�S���]��bb*Nq�-�,Nrh�5%�P��(-T�~K��gi�[��MY+���?SҲ���y}k��R�e�`��W��2��6L���d8x��vRtb׶���}�80PÒiO(4���p�%şY'qQ����b�<d���"��\N��]�/eB����c���L�ʂ�i�Lk��b�r���[O�Z��:�Z��q.��ʍ�E*&��cam?XD_�7�0�k�%�����QYTX2���	�8&I��Mh#�O��l���
	E��&�ڧ���|2����bL�q���b��⚃@9���m�k/�����H{�/_�����1����72���s�ߜ�K���]�^ɈY!�
��Pp5vO��i�����n�(24?��æ��`t8b"LHV��f1�������phܵ>���l?���͗Mc�qM=�,��lW����F��zH�$��&�Xk��Ehu�xK]�{z[��kGB�&k
_L����86��Q\ʿ���L�E+e��<���GX��#af	�e����>�ɰs�B�-�@h,3�N����	�=���we���.?A�����N��YWn�t�B��/����~��jҫ�[}��69�j�r���שǦ���q�1��7�+��|��R��t1��Q�����2����V@Qi,��?:9RǡQf�0k��K��e;t�^-�U}����?Z/����h��֘��>S/��̓">z��[�Pɻ�yq������a���R'���vT[8�ΡD��{T�3OJg����M5���5$�+��P��q�O\Sȝ*����aA��;@��峭0�S%�s�5:���t��z�oo��m�ps��q������p�/�:�Vs	�6z_0��~�1vG�=�z
∂���⍂2�so�\e�*At�*�3�:3�Uئj��7��)5�!��.�৤9s�<6����2L,�ͱy=�rTG���/o�W��N$?R6ݹ�FY������.��#is	~�+h�I��]b(Q��5%ݔv��̥ͯ�$q��D���Q����$$��d�,G�$��W?%�x\���	�,���R���*��	������Us�HeY6աf^j/�<�B�x��D�)�-�w�ʝ|��~+�]-���{4���������GP��Qil��D~���g++Yn݉DF-{�o<���b>xW@�����ڬ���\X��:Kd�����庇��5z�e_:W��vm/H��C�1K� �����#֢���`��`�7�;�QG@�y(>v��Z��"CԵ�g�I�M�^	K���U�j��2�
b$�-\%`��ےv�U�l���ٍ'fr�wuN@ݾb�t�g���Z��*\p���hc��I$��0�}�0��j�*�*7;�o8U��Yf����#�P,f�9ְӳb���ݎA�Q-.��-Mi`5�m\0��������Ɗ|	 �Fj{4�1�r1��o�'4��Y;����%j�B�R�\�����Oڟ��O��Q5��@;��sa�/�7BZ�gׅ$��^+|�'o>�{s約3�(�,&����^�?�[�:��u�`�&� �ױ�kl��,!hM28Y�B�S�	:����	t���<���M�(�A�>Ȯg���A#�n���)�m ��!�šN��]̡���9yx�%�v-E&'N�ͥ	owڶ%� N�ڒ
-5�,�i�ۄ�իz�������bā���2Ya*��-�EWi���LTI�������pN�������(k�Y�}�{[�����>ž�,e��9R���q�;�"��O�rƜ@��a0�v&��pg����ǛY��Q2����Ʒ�xOd̦�&%7 �þ;hB�n���,��ő����9�>��2��ָ,Z����8we�;}Q"�0�O�F��p��PPX��h�`��T���E &� >֟�����ɰo�Tt��]�΅�St��iӥ�/�tL����uN?����<WAGܷ��L25JІ�����6#�O�nKi�q�����5ʼ�Σ��M-�W{"�u�?P��gO��=���+^0
�ϙ$�i\��1V�K� �L������c0~��	��8��\�Fˊ�P�G9d�]l���.Q�i�)�;�q������a�*��ÓiD��5�I����cԱ�2i��n+~�}�_bؿ�8�d�y�G���8̭��O5�	���	7��2;�E�1���f�(��yoWHC$��ϞW��;���tbqo�ݺ���.���������/04�1u����C��}.��]<�Nb�^��p:esG4�;Z���� ��`³Cb�^f�w�����7ݤ�pA��݉�	��������9\B��~��<�x�H�sMi꟥W �l�M�5�|䮵4��=������>�»c��:ϋ���4j�=���@��� �h������+��%��4"��JW��v��p��9%�\.kq�O�����4^�$Hcytn.��~S��D�p)�IF�0���k������G�j�*��&		�A�������U���-����Z�=<$S�Dr]��}b B�ɖ�?��e��J��Z���M��ӿvQ��jP��F�`�ˬ��A�\'�>�	�W21Q�ޣ��$*G*�?�,��"�w1�@J�0R8[a��%Q���D�[���{�/�%"��E��g"���`��.GR��gK�N=b8!�[�΋L��r�aSm�ͅ�.z�Kht1�[�~�coe�Mi����ʷ=�A�܏a��8�9��T��I7l/�kg�y�D7�/��
L�x%v�=�%�ڿS�A��nMG�%�[_��G���kXl$Ǝ�[����]�h�_��m��L����!�\��ʃ�q�'�-N�S��G�U튥:|#��pz�c������s���Li����o��Q%�t��N�"ɶ��./S?�ݕC=��sZ�Y� �!���w�}!��t{�?�-T��.�i7D+����X6Y(.�f�Yk�$;���N�������J�kL����'<�R~ߜ3���ZwC~�p���?��3����Tp3�"�������P�b��\TƉ&p�[�o7oA��1���ZM��Tb���[���/�_�KR�C�n�瑹}Gkc�Y�"�WL�s��PM����рU���=M���U��;���r���/��d�a$.��$6��Z���a�}2��g6�dn7���M�ʰ��#R��ݗ���jO��H�Q5�l��Y;nԙw{b�n��+��Y'H�ND]F�X�K��poYۢ�8=-��6�S@�N<�6��m�ǼAz��|^��h\�0�-�fO�v�p�id�	�Z%�j򲠻�����p̱Ĩ)\x6�mo��L��7�Ÿ���̛7k\�\�b�z���;��Q\N�Z):���p�%�j$�3	�� H�~ �K=
ʯ���'�s�Z���i���l"�������B��G�B;&r���2�������N����,�r!PA��c� w�5��8HC�pl��&���^���q��0x�%S��⊱��#�O��C�xW<������
��.i"���a��7[�����TG����a �"����Rb�o����q�go _� R��F3
~NΖ��V�!�2��ܭ?�l�)1"�/4D������af��?3��w�2��Y�����9��X
�6�\�D�>�5�f�e��Ơ��t�z���f�v��t���P�'�8k���.ݳd?m??�5���``@��0R�-����F��Wùb:�Z��S)c�Qۊ����|`P9l�	�2���p|Y � 4E�-�T��g8N�ʒ0��Z�|S��!�j�n�l^�V�8�Ŋ�:W޹�?Md��x�P��h>�ƹ���~�K]3;%�AJ-;���l4���|ר):�d����KW�(k�ہ���z��Ɓj���� ��	=��>Q��6"��AtdyTU�a��3^���{l�s&��d<�Q����f�Q�HyV0^�LLϰ�U y�y��*������4Q������4�:Hpjv`m^�}�k����`�U��7�[�������HJ_-��oi�����f��$x0Q��dbp��S�>�� /�8m�m�o���_$��(�穖�P��.1�c>?;w�~��4A�n���Ha8SI:G�S���Q�i���Q�'��d�'��s�� CAf�ZO�:��qf�tJ�殎���y����y�|��f��8b�yߪ��=�{FIk>?��qθ�x6��w*1�xN)ŋ�2�-�5�����C���s��[����arg�͎!�$6m���i���{���4���G`�_m��{���V����J�"Gj�n(��j�3XQɢ@딞P�s�����t�}�(m��6���V�Չ����lJodq;XY�u��dL�����V���t-�kMܡT|vC�؈ �#Ƞ�~�'�ĩ�(�jO�(�k4/k��|UI��EgMۦe�5�m�_�j$�B� ��l�Ξ{�
ל�W��j}m��	J��3�(XS���!Z�`��D���V�N��۲���e�彈l�b�Ew��4��͏�U��`��^�++w�\��pE��k�Z_�8<���9�t�hH��8�[f+M�*x~���	�z�����F���k�*�~��S�e�9 ?�K������!��w��^L	�y�t25��k�H+X���*�Eu裚� �fd���ߵkCBl�I�#�4������R�r�s��.�����ݼ��#�w��90��Ѵ �����'�x׈�bZp�)Z�ua�����Y��e��ɳ7�z�Rn0kN���1
���Or�8T���NV�E��	��l��b:}+)c��bk���M�W��,�h��R|��6�C�l���}(9��m�Q@����X�;ĵ KYVo�W��uv�ώ,Ը��&}w|)	�,�ݤ>,��M��p���7�c��S�+	�RH�3�d����c��Z�Fc�Eܝ�p�Q�.cB�0gI8TΒ'���`���ď��#E�(YV�q,�?4��v7�" ����zr��⎨c�`7�B���`�J�hۋ\F_;*OVu-��:�#�[�腀$[�9w���,#K�ξ���z".��nw8�z+=lX���%+�r��K�8��=�ǟy�&��â8����+�����+�/]THΕ((��Rk�<�^ܺ�������{D�?��<�)j�J�w�kP�W`D��/͓��bQ�Hg��6�.[J�[3/>�@��2U/������-����M��'�il��3uri1�k��� -�3k�a���_�c�>_��{~L�gr{������h`�%�%��{�ɇ]y[<�GJLk�AN V��~.�*���z r�)B�KmوR���2Gқ�T�x���=zz�q�G����g
d����L��պ�mc5�="B��P�J�*q�^w� 9�0������sW��h�Z:�eٕ*�	*)�}��*�q�1��� ���o�v%�����D��i��\D?/S >�a1�`\Py����􏰕��A���s]EP�qܧ��\�Wu�f�yߣpނ�X��I��$�@v�:���'�E#c���,J�YpG�c�����gk����f%�07���3"���4�DE=���;�}��Bb9�����j�.�������ٷ�ݜ~zUɛ�ֽ��+�Y�x�
�?q!���	��e��5L{.Ү�7�z>��lF:��(墇��1����a�	�;X����J�ܥ��oҎ4<v -��'Ʒ}�`x�k<�a��2<�f;'���)PT�
T9	��?�c��A_�J���.�T�Y�-!mzyO��N�q�]����i�/rn�_Ƴ1��s�-R�8���x�Z�S�����7V�V��0��49~��)�U��|��+��J�`ǩ�
w�J�iM�^p�j���3��l�YuU�K=?I�X�4��8K4�S!���rh�fz��D�N�u�˲ނs�˞�M4F!��Џ�MѩC�Ő�A�x�g	�Ea�2יz���^B�#�x`�.����&���!�q��~}+O�9%`��T1lCy0�8��QM���H�ӷ�G��C��	�������jS��zA�Q؃��yj�b�H�$��:�>4=��"�M��+�7u��Й%r4�m|>�2{���y<�����G{zs�!�5�gc�����E���A��N�$ŧJ1I�q�"�ާ͢F����I�r��x�68�Ee,�?r-�\8߱��p[ 1N��5)��?s�%�{ȧ���F����F�ΩS��1G���+	'���l�I��A<�?�:GE�
�P�w�rW(�����%I��؂u6��L��,-g��0̐���Fp�?���i�+l�u�J��x���(
�*�Bıy*P2O$�c�V�N�r�^��7�R�!���8��ݱ�bʩ����#���I�@ầ�aK����/�,@P��N�hg��AC�-ٴ�$��BtjS+08���TǾ���g4���zQ�,�o��v*ܐ�be��N��/l�/7�>�@L|l�Ջ��ؘ�;�Da.�� ��~��^y�6��'�
�KpP�
8�T��������Z����b\�=�<J'H(]��m������S��}��8
��$�L�<zт��k5�x�`��v�=���/�2,q���g��c���#�.�8rY��M/r�+(��h&���٘�Vc���9Êf�n���wP�`R�N'Mw��s��t�YT{)6��f�C]�q�L/  	��ϻ�W�s��U�e������֍=�͈�^���Wy���>P��xf�+�l+E��J�F,�6�,z��-=��A`��@5S���GM5R5ĪBt̓R�(�����k�
�RpHU�N��p>z���Lsž�#�ԓ�F��mG�(��߾��
7�7�I���3�Ҿ�o$��Q \��s���,s�'��=��:�B��W^�[�Õ�XW�%o��(�<�xu��l�>p�UN6���i�6��<�뼐p*��)��ra�(ڡOP$/�����ӽ3g0!����X�=����*VLV�6��,;0�.X'�NO�u�w�?�{����L�v�h{��g���6G��t����51%�Aևd�|"�/�.��$5�p���R[\����[��o3ܱ���3���R^�n��t�C�E-'�A�,_e h�Z�z�&�U#!6�����O]�i#NO
ר�x����(�3�&zo�_�u[bq��ޞK��l��	����	�J�LK4)�b�D�M9��!q�`�Ъ��6tLh+�?M������֮�X���du�]�bF�pL~���쨖��f�i�rY���c"�È̄<���m���%<�wxXH.5۞u�"�d��[�y$4��=(�r,�\�:��Z��O�T����'a�<P�W_���� �;��'pmI�\�&PϪ�ѓdf�e>�iK�e9�đc�)�����I�'l=��rH��U�|XlxV64EB    fa00    1320�_`m��8}��`�����e� �B��+C#?���ڜ�j�E��l���J��cӶEG]�D���t�[�O��}�Fz��a��Op�O�$���*'O�e��[T+�.F��>��95��WB�w�e�t=i��*�&<��M"�'�^�����9?fIx� "@���N�F�<��:D�#aC������ ��/�(W�H�v�,�"��5�DzgZq�^E*/mFFO"����H/>�s"�7��}8f���a��1ja�KG4رW�Os���(��i� ʹ�bٿ(Z�����4��u���0��H��t��I3���Cm�+�!~ g��1�����֨	k���y`6M��SH"��u�>N�x���1�
�-9?�wj�g����@��y2��X:�G__}���YE��\����; S��ZP���Љ�G//��e��ǩ�R��&(

�x�RNJ�eAf
�����Q쾤,�%tca�2��tV�|b��|��Q�J`d벨�pZ��#cz���l1�# us�5�h��?�:����#���9�Z[��k	|%�)�[���� 9C��ؗZN�!k�E��,k�m#д�AbG�*���\>]�5���T5L!��撡��S�P!B�kHE�9���z.����&�bF�3��&��Hޓ�x�U=!�	��X�"z�V�Ɲy��������u_P�P�K��\Fu�zb��8����mt`�{��1)N4	!�ϱ�Tῄ�tk`e:�=���Kz��Bn�O�}�����a,�A$)�4Y�� �4�]��PH���V���T�E��:���?�����˂��
�������)7=?�遻6�T(�]xк��=���������-��p@3�H R�!B?G��_��\��@��)��<�Zډ�rg$�9��#mi{x�+��.dbX!���2����'/���>h$1��畬��F�KJjK\������&*�*����{n��˂T��,^ٷ����e���s���	��l��V#�5BB�	��ٶ��t��F5��;�!����'ՙRN���T�l�W�@�*��Jo�S:�8��n�Q/ù�&��.�:I3'bG�/yģ7�ȊC����Oޒ&����󽿺u��χ��P0�Na�����b�����6��V�\�Vh�yRchΝ��[ ��-E~ =e�*�;|�z��㥏���9��l�ʂq�w}+�~C)�W�L�?��"�:�����۴�t��yn4�j�J�s��)%F6PUl�^����ls� Q%�/_��7�B�U�a9Q.��c�W>�c�x�>X��;�}�č{2��[��N6:[t:��lh<��Z��K#�	�����;���B�ݩ�=�/�0e�b
ʳz��I
������:��|�	;T�n�%�{
������:2>��Q��`��	��$1O/�" ��X�%Xg>�iy��ps����^�l�l����.%[��,�~��y�2v�p4�)�m�����&�[�-���pl�%?�����B�K,�4G�B�Pߒ������ZS�\#��\P�K1,_����Xt�V�_θ��F�(�B��k	i����*��
X�8k�7�6�ƹ!�V�K^B�"ߊđ�uI��2�"/v3U�U8F�h¼1�y �=����Ŋ��%�bE�Hl_1y8�7 8d�C�DR�<-g��%���|�*������ JБ@e0L5R'�ٍ�CECxHB��hUg���r"��;[�����޻\�u�.fܹ�!Y�w��d8��1'(,�q�i!ו���z�s�#]͖ۤ.
iP�`!l���d�M+GӾrCYE��1.
��4w�һ)��DlYI�LO	p1&�'���@�a�|� EPb,���u�_�fR��A��zq�^Fuc�]v՛��U��(��ºk5q��9u�C��z�K!?I�e��#4�&�Y9˸
��p�S����f�'zR�}(���2O�f��(��v�)����ɲEC�w̱g��PM<Ob('Ϻ��h/�w��I��l����g��vv�.sAXחȪ��!tǱ �˖�߆���?"6$xW�%z�QLq���L(,	�������6v6���Q�vAv��!p������I�5{�X����⍾�|�	����R3�B����k&Q~�E�` �Fۥ� $	6)�~�����F��ւ,A#�K�+4(9�@���P�~�'��I�n��&Z�25MW�?�3b_d'���=֢|�[Ήu��-1�ü|�a�(z5��z,�v9�5C��('x��y�:IAO�.�����6��<����Y�nbOԆ��r�[�U�D��
��+�=[��f}JŨd[==%��7y~����em��;&x?.^��X��L3,��{���>�J�*`<��"EA�L �����A�h'S�+Ҙ#����3[�?
�:)bjK&wUB�i�s�<�%U�M��J����+ ��ҙ�]�f*�T:��8�����QAӏ���H������R�j��\�`�ν*��&*ik�g>�l|s�W��S�w8�_�)��,I�/Y?��c��+�a�Æ�0�,��.W8�Ԭ-u��EQ����>C{_yq=De-��g`A����*o���ٷ�g.TQ��Fzi�@g�aΒ��ͳ�&��I�5f��P�i�x�q)��zi��B�d�I�c �w�D���5`��\�kb�VT���YhbT���8��o���6h����'M��z+�X�\���;�-�eOq^���>:��2 ��~/z��N��cZ^���q�uR�듌�vj�θ׊���C��	&������K���p���i��z�t�.?���_!��:%�AD!5G�f��	�D:H�ds���_�W�!N6b5z.�j�]IP;��#���aW%:I|9��"r�����'��,�a�BPt���p��	4��ąE��7���oȡ���� �?��=� %R u�F���y@y�O�%��QV��p}�	�q�z����G/ �o�=ܼ��W\��Y?�7������P��#���g�#Wf`�`:p��7���Vk��z�� ����*t6j���6����m�(9�W�ǎ��@\��k��2�������ϛ�!Q�y��"�����$�6��/9�[kK�j��	h����n�l�X�5{�W���-�����h���gP�/!�`��];�����8��=r����`:.d�����/�|��H=U*�!���<�dw	)����1�Vᘉ$8�o���:u��1��I����cwAN����|��Ãy,�Mn7���Z��4`��W�h����а��ڂJ���5/C�1�t��u����&��� ʧ�J�-�6����К��sO����v"�Z���fb踑Ax~�W���gn���z8��źs��������=6Nb�~ ���fڇb���A�N���ga�JuA�i�{�w:<���~	{�[�~��IXY|'�ky���,�o+��8
G��s��x$y�I��n��1���]���m��C�=)�D��TZ�9�I���>3E5�z߮���gb	\�'��������^F��͉�wr��G��N`U��}k�1���Y�ִ1��T{���1��F�xw&��H���5���ϔ����׉%��m��@d��V�U ���Z�JMΎ׉��V*���X��`�tg(��A���i�p��IjA]�KկW#����斓hP*���P�����Ѽaٙ���M`c"����`~ʰB��qeM����ٰ��T1h�"
�Zq�z^�^.�^�?v�7j���y��š�j�u
���S��Ș�E����T4���������x����#�0Q��Lz
ʶ�-���B����-^#D!�#�1q�����;�&��;RN��tΫe8�K4�~���c�e��i��=p���} �G����6�g�+C]��f.<n����9m�7�#��0f,���,	X���n|��N��j�`�I�u6ʜ�]}Q���gs�y��'�r+�����rp���dI�>��S4�B��a��%�\o�#x!~�����nA�SEހ�g��ɮ��d;�N�6�D+�����g�)�vu�m�L�t.>��<�BJkɏlZbS�"�1���V������aZ���ϩ�ًy�B�N��`;�:��$���AKՒ�#��a��b8���D��ủ��`y�=��S|�u��7�`K �y�DU���N��@aY<��9Jݷ_�z�Sx��{-�%�^��Ɩȃư�t��8�ab�X��sAtNOB��|A�2
��֌�Q1h��d��iA:�0�P� I����T�E��*7>mS?�VN)Ś����/����I0 ��z
�&�J�W���D��v��F�]M$0Z�o����y�8��A�#v4��4�o�n��A�������<��>?R��;�����y����[�>�Px��f-�
uWy�0���������ٲ�=¯U�_J���
+}�U~�	�E���Cσ���y�w��6�ASa�cw,�ъ�ζ^p���eb:7<��l��Н�����e�E��\���L%��j5^m%hQuzv���.��"!�*�R�`�#6*�d/�<V��
��l�	N��KGg�`�'_2ﴰ9-�t�mG�k�����X���yBl��%��ҷ|��%WvY�:���tw&�e�J)��p�C����	���
�G����N=�'�(q��n~����C����W7m�	߳���g�_N�21 �QP�nT�#�B8t�A��f�V#�}o-'am o���'1�H7�!B�n�.�o~�,xN��+�W����)XlxV64EB    108a     3f0�,js��eAV�>���f(Y�Y��#u/x�/ �*��k����`�`�E?;�+\U�F��s�q�́�!��2NGs(�yu������bծ0El��뀾rQ���'?Sop�#��>�ŐT��=��M�1dQ��|ɟ��8�P����&+�6�����{��f��Ƞ�(C%�Ö��	
u���	�D�.���ݡ��YmBMb���������������Tvud-�:Ɏ%n �0DXC�7"�Ǒ�պ�M;�Gq����F{ݟ^��i������	yM �ٜ!Q�e��w (+t��<�\E�W}'�[<kB����f�rM��B- -!�!��Q��z�$A��������H�.��a2Rh����N8������<�R���C�@aa�Ŗz���P`X�i|p�eV��mvJ���jj��&�g�ޫ�D.b��g���L�
Ժ�Ōps��K�_Y��%V���Q��V�-mJ�����¬w�P��+/|�"3�����l�%Lk~�ȡ��mK'"�2T����0*�@.���QJ�k�����m<��������&�m�m���pC!��r�.q/�>���y`��:�.j4Q�Ĭn�+�V+���n{>�{���%%��/�8=����#�(wEKS�|�t
5�h�X���8>�P���V��rn�f�����a�Z��a;Ur}����m�aF ���0VB�v[�@�8�
�筙�B�Ĳ����%{{�Z� @L���V<�T騻IlD�lmtFb��ܖ��It����p�,��9LV�uQ���ٙ<A"B���{(,��e���RF�&��\�2�4�� E� gɂِ����n��,#߀�꿿��N��7�m�G��y7.�hkݔ ~X�y���j�Q�p��1%l��S�,� M� �#\�s��=do_��iى��R����_MSw���*{�+ �R8�|����_�db�UG��(��74�]���