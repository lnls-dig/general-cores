XlxV64EB    516c    1020����?6�"�Ac� <�	�+)�e�	.���pҧ����S��?\H�"�����;�yk��I�h~���ܮ�/c�$t���wqe � oɺ�lQ�=��<�3*D���2vz����zV1t��pDc����y��1��`ó	� r�5��?���{~���卶�7�/s�,��"������4�j��,��
y����ĭ��H�Y�vZv�Ϊ��&U �0����!�T��\�W���:W�;q	�٩痗��AN��J D��Rp��.1@,�U����Ԟ4vq�E�w�r���(뮦}�6��`��Pb�&b�*��85I��uPp⽗�����c��� S��(�?ѩ���^T��	�_�]�*��lS[��Ş��/1���%_@�;�gR�h_�zl���s���"�m#'t�Ԓ��I�\*-=�f��٪�;�>N�g�f�Ђ+�x�>y�Z*�\GTS��V��P�0AƢ>���9>­P����jo��@\�'%�\xW3��(��议+�x*{��:����j3�ŏLi=�&�P����v�Ua�ß�g���Yj�P���9�k-�����A�_�Θ�Ai��9d�o���ƃe��,*��8�VQ9R����Dj��o��ײӿ���	T�xS��P���0b9�B�H�ĩ
!�&����z"�W3>��z\����ju�و�r����l�����4;�ת��
LWt1�~u��պ^��o��?Q(�A��h\��.�ͬ���BRs˾�d�6���kP�6:�����p�@��0 ��A��<g՘m�m�h�E��6��X6�,m�<7����z6z��Wt��Q�a�wf�@����������N��ir��¹^�'�����f3�����֘�79�BYڅ�|N��5�MW���!����#A�7WO@�"[�f����4�#XK���� ��]���9A�.��jl{�O�h�育��9��y| `MOA��a���
7�UC�l�J1*d�3���BX�;�.a���vع�����Jt���!pa���j��'�������'B���]��(��,p5��8G/p3I�#�0��Z,���60b(�e��[�.C��K��+�2)E��DO�k+�I�ֻ��o�R�3��Q�n>|�|[,*��fG�����(���e�'/� [��EL����_�-}~Ѳ�1�_2����~v��ۀ�4�,Ӏ]�{���L����d|�m�������Ԥ��Eq������%��y��m�uR��ä5����|����U+"��u�@Lx�����
����sg;4�5�>c�6�#���;h�{�S� ��u�6�]��	]���!ư�&���?�<����}���)�X�8_*eN>5�)!�l�!�\�Y�[����)�����o;���v��	{�*��<��$��+U���������S(v�Ӕ�j)q�`(�*��0Y�.av��R�t�į2E�0�i:zh�֓ڮ�����h���,Q����_C���n��@f�gU)���c1����
����0����U�_�t�ib�� $���
	���I�:�\����td�MQ�צG�2�* ~q;�����Z"'C7d!]vAY��k�
[-~[p��r7,��X�lQ�Q�и]j_k	.^�R� Ŀ3�9��ӷ��=L��b?"�����Ul-G�6��Z'�qt0-35�ϩ�tˉ�n`!�g@Q�r�j]�9:�)Z'��B����{��,`x&�������uJ�j��V{��±�Fv�{-5<��mf�2�6i����P��}��(��rĨ��k�5�"���S�:F�32rX������қ1)[�*��k���d{Y\i�2�z1�+4�߅1w�τg�Ίo��|�˥�<e�&YT�I5{���bb?p��6���4u*�0�#7��Wvk���O$�z��� ���ᣒk�4������?9�uS��Y�E��3������کSH(�-۰|�fI\]I0��@
&x�f}��-{���Q���a2���Uo}�m�}˙Q�����u="�Sv^� �+�����UX���(d�8�+53�~LW���{r b��j�F��7т�P��ν�U�O&��b$�|�<�e�	�LVID���0���k5Ij��G�ă|o��&^�.߻+�m��6�wY�b"j��|���s^=T�x����k�,��P��)r6�E}��pkM�!��R���z#�E��w�!�AK�ь��
�����hl�M�u��z�.Ϣƞ�]!/~�'�N�RC�c�4,*։t����sm�0\�Es��D�JAqn��e�r���O��6����Qg�!�Y��V?%���2QOB��@���83�ٰ�\*뭩=���������_Eey`E�Y���}@q]+q�5�ZU0��f܅�<=EZ��8��_!�-��V.��d��Ky9�c8���$��t\/M���b�@8_aդR��R��]�b��!�#��Z	�8?0d��w�E5�p�J:��̠�6��������^�^�Z��04S�@N{�����{��r�܂�l���j��Æ�B8�bƗ���Ac�����a��1)����|��Y�CQ\�F��(y��Ǧό����5�b����:�nɭ���������ˌ�A���uB�Bb���f�:���:�jK�{�T�5�k#��t�}�S��tC�O�^򵈭kL=NA.�U;�ev]k�D��w��K@�ZU�p1,]���z�H�&���$I4�۷6�%@����q(9O���@�c�q�ӃR]UW�YuS��%��؂5WE�Ã7�/U� �q��<D�q�(̚����F8�O�ז-ih�N�'T�Vr)!�:������O��M��ZWFz�Gb�ţ�^��Ҍ1�}6��(vs�x"�4�0�W�_�����> ��S	_�LA�����\^[�~�
��倪<f���Q�3rp���by�|���C��)��zx�[�K��ߴ����R�`�����/*��=��a��j�	��JM�J4B���ǰtX��t������~F�$H�,������7��)���}n1^Z�h햑�BM�-d�][ٶ� �/1a�H����g��i� :T��]�����i�6��q������)�tį4㨙<��1�B$g[SP���-�|=��v��O�j.��&¦��n��P�	�,#�Vk��7Y�r�{�fR�}�!�t�?r���l��a��sx���[%6�Ug��[w�d�`�� P�"��(g��]RH�AW`�g�=���yy>����>F��Q��P���k�]K�<O����ء'I�:d���|$U���{_qt$�oiCX	4�����M��2�I�!P׉63	�1��fr��`��j�oWEضt���n*H���|c:��$.vD�z�*��z��&�h6َH�h�tB�?k�A'�b놿��V�)Ԑ�
eU:���4��>������M��S�����3���a�<�Z�+<���
Y��D��������#Ş�Х���_0�B�0�{�,H�gW׏^c=�|?n��+�M}O8��� ^�7��1J����yeat�%�'Ei1��j� :&�K���\'�f�O�O��M��{��Ze���`�E%��ʕ���X	�!��uI�s;x@x��'���}F@~�e�,=fo�����:��I5�QY�WͰ}�*�'�����
Zu(H�"��T�{������Z�R�f��F�o
��fr�L�g�-���W�/��'~�[�-�`�����0�(�̀���R������g�\|���@R��JD57�����J�Wu��yw��� ���r�.V����`PO�����+AI���Ŭ�k���mw����M+��y ��2��@��=�iM	�Bإ��V8aQ#Yh:A�u`��
�6Ҥ�fh>Ր�g��|���B\�����SZ'(G�:ḇ�f=9l?%�R��Oj�:0�J�6�8����E*�-7��>İ���� ,|�8=�QKF�+}NT"�Q�������8%m_�I��x���s��%��L�${��n�i7t!`�P������-���E��A�V���ޟ&