XlxV64EB    274f     b70v��&4��u?[W�����5�����|hXS�hKC5��rqx>���r\)�٧�`��J߀�B�d��@�����Y�-2\���M�`��96[��^��O�.8�'���4k�cQ����'�Z�v7�ڠc�:�)����,T����&,���N�������6����/���JWm�k�V�g�2+Εk�����Ǥ��ƻ�.�ĥ��7B �Lg١�"Ya�Im�,noۥ��ֹ.fP�-|ǵM��O:��
G����߯�5���\ �7����_����0\k��>��:��ʈ}�X�x 2��Z�����<���t#MɛJwON�ػ\����V���ۋ*_�XP�cօ��Ч��������Aq�Ԅ��5�tJC�:��D��I*�S�]��ؾO�f��6Z�۔�_b����w[#��,�:$v3�����[%qK0K����"��.�`��I�@�P�d��i�0�/!{9�!��B��P�	G%�+�,�HbǏb�O<��u8#(h��d��h��z17�,��BvE��d��*���.��Vb��ăP�;���d��A0<gn5��Z��a���Ф��[sGd)xU;4f�9�3r\��>DbW�>U�訁��p26�D���É�/�^8�3���}'�㕪n����܈��f����<��:T��K�\�M�}��Z��g�j�τ�x#��$r���!�/���-q2�
m��C��C :Hͣ��U��$������o L�
���OP6>�HI10�������g˗�{��_)��W��N��2�$ܘH�"�]Cz0�H	�q�rf\7�z�	�����>��c�)M�$bi�a~>��޻n�EIg��>Rs���n��琊e�	��؂��BBǆg@�G�'����Ė�'��24��)P��Z�����̈́�r{��Y67cH��X޳��tqo�"���v���?q !���[;�Ԋ�ާ]j�A��cU-����BCp��&�D�V�f}��Ҍ����M��ݨ����;�㺒���HS�j��gA���3EŠ�ut���M21�0<�#�I���!o%�b���Ə�y�ߔ	~rn����/�W]�@��|tJ�~��{����:��!�Cm�c���1ڈô�~��:,7�,1�"{q{�f��e��aT)�Ύ��?��}��3(W8J"i�ߕW&'��p.泋��$8� �'2��N�F��hF�M*�޽��Zk��Q�a��bj��c�Ý��%$���3��n#����C���W�O@���7�䂫V�� �}�XH٫�n�J�G��r^��,ZUг���	����B��;L�����a��(��}ۥb����H��Q�#}616���T�����ν����u�RN�FV��
�M��C�=�w^�p�,��?���܃������7?+Ѫ�o0*+��	O]kX�+��>_8kn����~�L�"U��Z�O��8h�!q�3E���+��.��fٟS�1���<����9*H�\\��ly�E|�<�CwR�a��D;��X�}��:	�SR��߭2�7p�=�r�?q'e��>��j>��d�MS�⅙��p��? �od��!���P����a��Y�Mx��P�@����%U��|��q�	�3~�ne��	L����^��h�b�dk����g�wU��.4
~7f+�Tu����':�\O�KH�hk���f�T%A-R�V��0�8���z:.?��G+RP�^сPQ��F�dH0��cv"q]�>I�䜸�	���}�w��]��+��-RQ�o��o��%�u�Dn}��m�~�u �l\oG���U}��B�MHK����l)A��C��Y�BX
`HkX��g�Z����F��bT�m��lM ֚��$��$.ñ������/��*l�J$��y��3���B���`����v���!,����s�u��AL�R�~�nj^W��AHcڡ�w�`ԝ�QϚ��Xޗzy�����o����9��߮-�t�$�d98EOTL��������Q8y�R�Uu������j�����LKwS�w�D{L�噢�����ȱp;�y��G�kG�� ֳ�(�������a����ןO7�/�����H!�X��&d�En1��^�Nl����nU�0��Uuz��ǌv�p�C!���D�Q�j������
r�nˠP�Z����qnp�e�Z�R�<&���+��a�C'j{�A�^/a��M�6P��}� �����ng�e����b�<nH��v�����y=_L�+�)Ѳ��fV���Lr��)���/�;��oa�)���� ��h:C�l�;��#n�OĄy����T�B����yN�t.rg����z��!Z�)_�4�3�s�]'i,XUjJ�m �gY�J��Z�5C�qTA�ݸ��'/�i�~m���:�S�R�lTKMF	O����f��gX��2�>z��F��<+��"5�'��?������Vp`9D����J�=N�B�\�a��������NӰ��*=3^��!(�i���YTy��4�/x����gs^��=�nЃ���0�X��*p� yU���$�@��疻b��ן��	�
�%t��֢�g�<����Ub��B7��^�𽟒�X�Kd��L��k�n��}���	v�%���Ϯ4�l�)p�^�W���& �F�}�*%���Qt5|��[�e��3�j=�W���y����uԗ${�����-k�У7���Y�/��&)���Z/�zOe]*�Ѩs�;9�����V�-���N�tF���_�I�WQƶ���ʬA�ө����i��!���.
��-��$��a�Jb {(S�=������w׊�g4