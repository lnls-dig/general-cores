XlxV64EB    3b8c    10502��Wn4����W��zH�:��b�6'�j7?��.�"��91���*(�8X�T���A�� ;�=�P�AG�-�*̞?e�aW����A1s�@����ܼ��f8��ѿ0-���C��/�R����_�|Wiu�����'�;'��;�j��[���P
;��,h�v�6D#	ʶ����zte�Rf��G��R���|`kh_KA�3$ڌ�@���	�c�G�Π/ x��?���l�]�F|���������AW1e���b����A�l'��r����)^ N�t�����| Lf���_�����)��d�k����ը�DIcv���Ye'���� 25�b�!Or8y�˞��Q���aO�9oA�DRd��܃aNB�-R�'ʷg2���W-�#Ӕ��2B&آ|d�ha�T֭�"�@��e�DT�U�.���R6h6��4�I}{rФ:�hg�,�J�i$���K�miHx�	K�E5��y����Ϧ��G;A��c>UL��|1i"���"��)S�H�>K�U�p(�9�R�Ef�����#/Lf�n�F�(B������\��2��e��f��6�cK�����"��N�1]kV$���D�:&��غ��r���g�P!�Z��N^��D�jw�&z�Ð�+I�ފ�n��$�)�ѝ[��B6 �#v�OtNC����z���ݪ&Ś�|��j�2F0�	I<�.mঠ��fI���hQޛ��oK��)Ws/�J�0[0\�Up~�n��U�n��Q
x�g�� _d��a��޼p&I�R�w�yXA� c w^��O�XPP
�y���H�7�A�B ��@"a!+�m��9��fkˇ<w�R�SvN��aL�v�C����c�.�Q�^H�p]?�7�t|����7�.A�L'��Au5R$c��7ci�jѠ���}x
d��.���}7ȯW&\S��´�!Q�vj�eRZ
r":`C�b�˴Zv�1�/��Yӆ�x[fb#�v��/j�i�������U{�Ƥ�?S�#���y��R�i��ZP�9#��*��n~5'8��������tĕ�/��~�=��c�Mz"<EՕSM'wY��Oy��nM�D_�@��~�!�Vr?!sSq��"��Ƥ@�������QK��U��[��2c���ƨqp�	�%#Gܼ�=+Ȳ-+��s���Z���n����@pD������U���O�~+���w�kZ�Yp����
fp~nU�5�eϜ4�g�
5�����^�Iq~��o+\^k�--t�ЅQ��FK��_��&s��b���Z�cV��_�q
���,�7��(Y�'H!m��p����8K�tB/����DJ͇��&0,�e���-��ir�����dE��m)4��;3��uʘ�h�������‫��a���:�f!=�u�ϰisV��x�y���]�g��v���d�ȰӬ�r���I���zs3V�ؒ.���`�2����O�\����I�zh������L���l��C��>�5i��b��M^�
F������,@���-.�K�B"���[����R��ڃ�4�]����0�0_g�o��=x�Z�-���1���m|�;�Փ�\�Q[��
;6h���X��֤67�5ݗ��xl\�	��ߒ�Ɩh���É�������*��H��H�a	p�'�Ud�	���E�2z����g�=�-�F$~X���'�;�9��H^�⢲Lճ��wu	e����������ú�:
�~$˒8hK}��7o�g����E��	���W�Vf�x���TZ��àt��Π�bfN�C�0Uu�%3Ol��)�n�T@v�d`K�Cq4���ÕŜ�'�(����;�.�x��1Kc�.���q�YE�Q~�B��f.$u��#�UZPᬽ	I��1�%�
+=�A̓� S����3{���H�d
�9�Y�݂�-_1�����b�;��A�e�X`Y���cY>*�ы����<����TC�����Y�V�z#F��~����j�V1&-t�n��jm�,f��h�E�2�Y�Nʤ/�$:�sQ�] ;�%A=<<�S�ZOH�H5�V�v���Sh�����]�y��gq,�u}�AW�_�"Cy"�ccc�A����Xf�*����6�J���}/ڴ��m���W���״�Md
�\u�����zs�e��P�M��!����+�8PAЫ8E���de��������I46�̠<(M��ݥ��跹�!A.�����ai�y\�o�/��P��N,�{���p��>"Ý��u1���[�	���?����#���v$d;
�c���]b�3� ����r�0}�nr����"QT�`�<eZ}�Bk\�7㯓�B�r�P[3=j��M7�l�w���������(��-R�#V��@�E[+"4Ű�*�X�K�[�!_~�&��
��A����d�'(si�A�'H���Sگ�ڸ |�8�V����
*��=��e떙
��8��K�x�h�������@-[�1�(4C�<[�hl3a���*@�e/�tV�	\����� �`ŕ
�.&IZ�������Ž���ҋ2+RN�L��G,
�.t �����<���~��F����O����&�Tj��!n^u氷Z�H�A$�h)~&��D�5K��r�К�b�&W�ؓj� 2���F��7TM��Jf�A���ɚ�f��vq�2��IU�`�Gĳs�W�*���N�fT=ض3њ�H�;�!I�L{JŤ*��;I<mE��~Go��T��[)83(h�l���YF�
��*&m���i�-��y(�!>�X�r;�i��t�	Y�[C������W�V��;�w6���e"/�Q��xn,~Lm׏&�b�8,M\����V�O=�b6뢖:*ѯ
�A������x�-uF�Lz]i`����,���i�(�P���M�I�	< ��n%I�=��6�}�2�?.Oٮ��8NS��ӎKU�Y�6:�p�fAbD�=)�FVm�Gc��v�Ea]�Lq����l=M�9�����AI�又Z�s���s㸱�-f�������o�tV� ���5 �塐1�o�����ʡ�%݋ed�������"h�D*�Wn�v��(P-ᗮIG�|U=�+�w��9�-l$\����p��q�*�)�v���u�ħ�1�lz8l��iav�/l���wz��%䫽Y�y�3G�{��}���*bJ���)�����A�>�oȡr�Ё�'@��o��{|�S�4;3�HUi�w�g�Ė��emU��!�r������=@)��Hq3�$��w��|ϭ�:�n��	�?�?��� ��n&P��˳����C6w[$�fS���S@�).�������g�}���`�ޗH����.ٲ0�v����w\4%d�%�����B��j�y�zi�1$����;evG�&� �ɳ�A�|�?�s��VEaw������c񟘬��R�)4��5{̗@�?�'���=�'���Sߺ���a��^R�yԻW���O/���>Q����Ob���yϥI�)S�;*G��ĭ�-�ˣb��w���t��zl��Pj�&�@0��УDha��n2w��_�eG`Cz�ɲ� �*�L"��k�~g��F���Xd���w�t�SQ����7�-��*��do?��Q��`�
��H=+�f9I�ݧ�X���SsrW��
<U[��G���b�gL�(I���,��zgq64�`+�QU����x�HJ7�#g�<�^N(���C|�u������zG���	��9d|h��O}�㭧Z�Rj�"e*C��I^����t�>��i��g�GJ�	_��� ?H�wB~W�S�'o� hxje���Z�lD.a�m{�GH����a�d]�|������P�3���s���8Ng��`&/y�n�
��.Ęn��<ꨭ��u<�/���"�DM#FVϗqkZ����q]��h�t[`X���yR��x��q}���^l�@q_���K��6�Y
U��cq�G�R(���6�<H˥]q����`oRa�!�0m�ʏ�6~�-NB;T�54�4y�/�u	/�D@��:"-#�QWiSB�l��4,�2 ʝP%O1_���#f�}+��\B�ˣp\y]{)