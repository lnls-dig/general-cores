XlxV64EB    bdc9    1c20@��'�C��Ƈ���7��0���B�C9Ҭ�a���<�x�϶�ł�%��d�\;�9�:�!�Wc8�&nx���J���̆je9��C���X�;)N�v�h������>k���ma��#9����j�i�B�ڈ�]�.9��xm��X�����{��O��	��P�}W#"e޼R�D��l����`�ĭ]d���E�)�v��723{��0�
�R��'�ɞ�O��5��!�`���%x�ށ����c�YCY��Z'���s�����6�?-aE�[3�J.�>�U�+0��;+����C qAzW��$�h�t�MHjE�Q�7���T�7c:�����}'yW�\^8�@n>��h
��Z�����A���i����̈́�V�b��Bor��	��A��*Ҩ����9����X~�JL8�2��E���o��3��V��A�����m��fE�Y ���Am�_���S+�W�V���ù>����F��'�ϊ��`?ڼ��vP\�Ga������[�jd+��?��~M8�U�I�s�7�3\�\��I�a�d��G5FX�Ο�*��Kîg���F	hxr�0U {V��\�.u-B�ˮւן^@�I1p�kM}��f�"c�����l9>s�1�@�R-��n�X�o؞��h����ĥ����2`��fJO*�`��>7q��T�OG������^������ȹ:E0W���Uh��_��t���݇����n�������bW�ՇQri���&w�kk7�էҵ���`wf�)�v�.��1�[���ъ�)���A��d����<������M$�;y��N��=���`���L�#���<VA��̒�X��<-G[0�t�)�k�^��&Ƚ���o>�')H��P�W��
Mf���ϓn[@#���Me����6�su����y�o��=nX9�^���Q�sz5��2<����x�N�%/��K�����&�X��l�{U������i�6Q�+z��&�,����Q��򑍪�l���{_�?C�Y]��6C�'0�Cϰ��C���6��#�����^$���>�*(GW��q
)ma��{�=H M���͢�SK��_t��,
��{E��E3iC�u*�b���aW[*�:M��r��}�ߟި��O1��"g#㱼�]�Чe �}/�3k�[�$jE�!v%s�n����Yl�`u	/|;�Cm�k���&�Mi^��(��J�h��g*����1�8��#���rP�@j�P%����[}��@�3"�t�NA��\���ه޹��ob{���B���+�5�'Z��66'a)F3�M����z�;؀����-6D���>�X��r�!��4�D�H<�e��:�:I�`D?5�Zh���������춆���u����e
(U_e��A%�Y �^��t>J-fB��kC��Y���k�h���{�ލ{5�{�����LT.�<�}��r8�yd�lb�6Ty~-<alM�{���0�I4-�R0��W����M��t��Kv�ĵP�xZ����^��|:�OU,̕+�L��j��'��pRD�I��@��	�*��)���*�t&�)�r����o��̖��D���I��s]��|�>�!`���Q��~�}A�H�E�����kD���Ȟ��
�6�:��Е	��Ԕ,��;�u�ZJ��ql,U�+�2�>hoJ\F����=)���w�d>��`��GؚUL�zB𯎬�FO6�����+;!�1@}�j�dX�x�+�M�6^�7Up[w�D S�-*�dcXD�+c��t��Nu,ZޮrD���Ob� g�wm�]Q�з��nʜq��l��`^�E�m�)uz�S�:d��H�s��۲�y��<mk�y���V�)�T��4�Sd�M�}��:����:��1�}��%��f�]4�\`�W�jgE��U<��K]wum�� ��9��S+'[8Ѱ��6����qg1���
]g��a�΃Y�Ւ�o�X���	���[��T�B��)�.zV3D�d�Uv�iu�.���Ytd
yN��	������8��!C������+91ۂ�X̗J$��v�>��_)��а���&��qn&B_U7z�^�G�G�n\�d-�I��[��dkG�{Y*���)^!�J���LJFa@OùzB-J�`��)�O�8�~P���u�ߤ|�Ə���[�e��Z]Q��"�/�6����rz��/�	��h(�Q�.2U	�ok�L�t�X-���'�R�; �$��k���˥�<��³�Y���d�68�5��C�m��AHt�%���D�A,>[�Qz%b�֌n�-��a�����-/r;"&(���`��HB�r�0r�[#ޅ4$��9�d����A� ���3�wG���O���;��:��g*<%pBఋ�-?e��ɑ��k?
Ab���1���i!�>~(V�:�R��ݠD���Ŧ��/Pɟ��f��Y;/�B���X8�"�~�5Qo˰\*�lJ�2M��g|��"���(S;���!!���:z�A�Y,4@�&��b�d0���WV����wx�Zꆜ���Z�/��_<�#�vw�y�����B��]��Tl��U-�ݲۛ�V�_����r�e�GZќ��u:���%pDD�j�v��GM��f�b��{�C
����n{5	v��T�S_(	��[��J}�0�ʍ�����f40������q!��z�F � q�!�b��Fӎ�< S-|}���	0��柨����8-�����ߣ���3W��$�� ��G╭�R�b�:�<(9����QA��8cbQ&�����m�e�yrӮ)&�o	,��cH��E�Ř������M[�C�&�� �*Nuv��	���h?�h��'Y�+i�_7OxM�z��6�p]%����dV�!]z%	0ι��(D0�
}��Z�[W�KcQp��g�W%�.�9�0i��T;nC'��n��tL�x���Ҕ��Y1�X^����::l�D���W�Y�k,xe�\I��y$�\"<�Ò�嶊�T��:R@�Y�퐏���AJX��e(�q^\�*�����"�'"����S.�0������d�C��)����k��53j�] �-\]�B�ݣ��:�a�O�Gڈc�j��CARȚ���./J��P)�Mg�٨Z��}����ݭ���K� &�V���@�ϑ6���GI�o���J�{���f��t�+�\6����v ���_�ܠ�q�r�Tn�� ��� S4k�U���;�aW�����x��G�H��y�nz�Gf�'
CHi�9���&u�� M�7]���syEv~c�R��cd��:E](I����O������P�8��h��$tCa�g� ��lyP[cL�,5�(��n��t{��
�E�q���u�ީ]��u�*�;�؊�,� �y�:�US�(Mv��~"������A����BLZ�����
������0��H�K����D�>�N�M"D����
ς�'Ǡtz�D({�@���Z�et~��Sf�Oz[���F�o}�H.�K��(q{�¢���K��<������.��E'b���.��KD,\��C���*�g|�J�|Ԑ(��c羉?V�n�I����
FV�#+�l0�3�k��� r�R�oA����U>tx�� ��r�T��9�`�a�q�';rO���y�*c�H����|�4��ܝ��>�C�V_iT k�[>�`rn�����x��y
/n�=�Ӫfx���XD�l��eq`ȏ�}��J��fŋZ_^)�s�����3�F�/��G5:���
��xA��=�3U;���eHu����5(O9-8�fg�z��x;Q��v�(aq� s��-�MJ/�	p���M�y|�ƹ�"x�X�(���V�(���9������Ew�J' �C��w	)�3���F~��`���f�95���:K�]�ad�y
i�H� s.|�r�i���� ���۠�2f@ê����s�]����y!4��</�!1%�P�ߤk�Q���9�wB'��{U�^2TA_��vF"L����/�Q��Q[<͡X@�P!���l�<��X��	�l'�+�h�' 5w���s.��Ov�^�_�2pz`V f'Gߝ.q#J,p� �0'�[<�۶>����?���1���s��o@�\ �f��Y�) }z��p������~ uq�p`�*�mr`�2�F���P��	@���=��Rw��O���,&���	ӓk 
�V�hQ��i-^�-#�.�S+ԋL�sL�A�?���;���sB�֛M#��3�g���?#K�mߦ��PW�C�Yx��T��+^�H�j�R�SbB���'X����9c����	[���?�;�Y����t7<�o�۴����v%�����3#������j�P�}�G�r����%��Pa��h~�j�*>�=΁=a;�0ۂ�8�x8�`G�����M�Hs�؃�i���}s%��!y��Y�\gѼS���E\�����ެ}��������r)�b�BY���4�ŅU�s/ߴK�x��.}n������?Q�U��Y;Г���R������_E��+iw2�:1��)47S��1���{TB�-,fׅV1� ���P*)M��AC�^�D\狃�8�������.�s�wy�CF�������ԅQR~<�\�Kv�UX�72B_#��$B�޺���Jp]w�x�N!%]%��:/��}K��:u���S�M�)��<��ܒH�?�� `F�_������9�(	��������T����($o�Tm��u	�z�r�p�{R}����#�)�]=�<
��x�G �;XeG�}mS)��Hi���#��d�J�����\��h��iZz��0�p��*��;�:��LBL�K�#S>�t����)��JZ��R��s
���WA?�����t�bƎ�_K���s|�$�[�y���X�8ST�v��������ve�"�+G7����5�M��W��u�������w��;�U����o��V��9��U�����7m�VP�S���E�=n�Q���ŝ�����{(�����ހx�Ļ~g����YUv}�H0/��@c(yܗ;����#��f�$�@" J�ݼ�X��K��k���#>� [��X+� �͡��i���}����Hi�e%��v�O%+5Ş�B>]V��ɍЙ#A��Iu%�h�%��o� fj�eQ�[.���_���.���z�~r9�8;m0��&O�s��W_xH��Lt�P� �X7k#�ߡv���u���-���[1�K��J�hb�J��Ѣ< �����I�H��jE;@|@�xa%ف��� �f�u�.,c�O��,�Ӗ��	��AwH��"8�J�	�CѮ-�0��?tT �z�HS��<+	��]��sǡ�M�?�� �'���][{�������$ǽJc����b[����B����6��y��9O	r΢�튏�e����R f�H�J.�ܢ�h wp�]�mq����*<�E.�oD�}e5\���P����)P���L�����K�����Z��;o5n�]Ř5ɼ�N��P�sV�v[�(�1����{��B���vC�A|�S�oɚL�x�k����r�5-Bdg]�u�&4���\�"�b9���oE��H�_#���#�z��y>������Wӫė6�S�1V�����W1�$�˷�%ts���	��a�:P�Yْ�Б{����4�$y�x?`��7%�r.��9�ᵘ�de�~Qpw<i�6�I�a�	��	rܞ�S������o��S�7Q7�� ����>�ȳ�5��J2����9�2=/[�/����:9�Cɡ��>�,�A��{~#�/'��������X"W�͞�.Ͽ]�1$$5̄�i.e%�ДWF/Tշ�P�n@O(*��.��P�ў�x�m��*�3�nJm��T��?o�ą�}3�"��x�)*���)�Qg�P���x�<��hW1���JH��0�� JuGM,F�׌	��:ԟq�Q�N��$���;��|����ss�U�;��ڐ�XY]��������F�>����:m��I�qW��S~_�)����U��e�H��e
��{@ֺ���D����Z�s��{ƍ�O�Yhr=��Rט٭��-Ԁԥ�z�XJ����L�{�b`���7��C�o�e��81�ɲ6�\����y���T�!�Q�WK�����n�&G�:�d�-����^n����%�-�u0�M �������8ǫJD!<ݕ�9�k�V|�G
���w��qJ^�^�ǘ�:��:�+��7�B�)yc��(��_۠h�;��9U�����n�]!.��i�g4���������25��vTX����+���$�C���G�]�Є�JSA���z��
u�;��������zQ���pRzH�0���%��]�����0ny(�,����9n�yw�KVY��P"!t��ڱa��^�yY���e��9��_��*x:��]��%�f�����
��b�:r����fo3NW �l�,-+�o3�A� �J�YFlo���c��*�TwI-HԠ�E�6��}>���zU�3O +���k�O����B���B�F�M�H�6��l�k�c��ͯ�nd>�X$���ȥ��E$��Ꚁ2���:b�1���۴��mkj���` �*b�D���[�<;��G�g2�~`�{<�Jb�T;@2�E@G)�1*O���q�����'I�;����®a�n�[����v"O*�*��d��{v�_�?3��<�T2���(LRp;ƍ��4V&눳S�^|�~�[E�2�&�qW��q��!۷K2(�B��J��Ƭf�&�ߢn�܌�b��rn	[p����mӧ�0V��y9�/��U�y�N~`/�9z�����V�x!����/�Y%�
9'�		�Tb�bd�x(�i�|f��'N#���X�9�?h��<��tN[J�u��uv1k���}ņ�5�#SM�x�*�g1��1k�����tJ ��@���m��uYsD�%.p5~��E/`����D��P_��շ�Ցq��F�����b���9����Η�!����T��^"+�JsҵN��n�ձ #/R�9