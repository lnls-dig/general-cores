XlxV64EB    8ae2    1a10�@�(���y���Z|$#��JW`��V��&6�O�9�? �H�������q�l�|p�|93�?�L�3�
�ԬMV�T���Vwd��L�y�P���� I��#Ol	̾X�ˮ�wN�K%�t��[������zĢK�͒��~Q͜���l1r}�I��ٺ��Yx�e��I��[fF������uQ�����8�H�L�RsS;�_3:��Y��=���َ[I�}j?�����'���j�v���+��D;x1s��D
�l�Ջ�����01~9�2P�,���ZΈMI��4��'.4󪩻LG+�����b0��f�����Yn���Q�k���2-mN[�`�߲�z����M��:�D��,#�S0	��wa���j������z�*���4�P��܀�	��A,M�:�%��{g+mxOx�I���Ku���	����A}��mE�b���5�*^�8����-�RF&I7;(�oO�,����$_���0����GD��� ��A�	I$�r��Ş���_ohc ��܍��sb�+�"��PgJ �
�xEG��}���3d&��w�v|��!��K�B���Pjt y'��&�D���`R��������Qa���!Y����?s`�w�+�q��X�[��3//}ʃW"�otͥy-�.ĺ���``A��1FL��RS����h�q�m��<O��3qa��"o��X,��_Y韫f^�V<sI�""���`C�z���T�;�t#s�<��Eq�q�x�ٛ� Ց�n��0�)�;��%���-OS襑������gpyu�NR�UE9�W푆�~��3n� 8���kѢ����n��O�Q��;�(G9��Q6�]L�9�-~C#�DL�?֜�E��O�Y�<ݖ��Iܳ�-l����5Ȇ���l>�����0hk�s��,��ϻU��ӈG^��<����V7�t��EHڽC���g��Hl�T�$��W���J�+��ʔ�Re7����ߍ��!:`¶H�Vt�k�4����h�r[�0F���o�M�f�-n����0�'��j��J+#Zi���c]'�.��ϴ�����[��`6��bo�;�E~�R��-U�g /?�/Y���L�~wͦI��J��d�l\�L�4�m�+���˺���3���8���NS�Z�S0��\��YW��K�4��N�6��F}�?�gq˰,��[��I�w��~���:9x6�Ӽ��$��I������g�TJ^����mb�L���沠�r�!e��)N�;�ή�Ǩ��Ҕ���;�MV�@�������o��_d�^��wђ�_�
����a��%��fuB� v��D�����X�:SE���d��b�D�w#� <P^�� ��É��`�Ky|�6��	̨/�v��1�t��U;�����|x���R�B<��=���3��D,j���K  ��tV O _or@È�t	�U��LG�T�i��'F�	�ݮ��-M����?��]��0���� *+����F"q:�����#2�f�h�(�˪涍ߠ���
./?��Fy
�W"h�t)��N��\{��9�O��DN�De�����T�i�6�[&�Y4CDr�t|�U
�cQ�wx)�Vq����$f�v��7壯iX>�2��y��2�X�T�>&�ߪ��f��Ա���,���/Mq��@o;��V�ؖ<��@�+d���X#�*R�T@4Lg�e0�ij?�lF=��t;F��)i8]�(��(� D{�����&7`e, ?b�#	P�c��A##�YD�k�R��G����2���[���3�y:U�kG�|)�Sh����f���u�a�Lcd��0��0e0���Z��vƢ�KMzXM�>�jABZ�`�+� z�%H��ߊ"��Y� ���V���Y�T@���6����;z��?i�g�e݆#
ǉ�IjX��t��M����x� ����2H-6s����A��������V�lW!�8ӿ�d��lA �PƊ���^D������h6���=v�h�&���Q3�)��Iz�������$'�D�y*�'m��zU������m7|�&�_��t�!� ����h �>��e���*
�6+�������=�wo�D'�� V1G��_��+�Fw(��R鷊7�r��	���P����ꍑ�ƨ�W�!��^d�Z*��{��.�m�$ǹF��z5�6�M��v�p���Lv�33�������JT�q��b�I7�� \c���S���Ze���W�K?	��X��{�<^H�<r��n˳�ʕ���C��K��S����b];�<�)�v�qu;����_�����F�ªz�ό�@���zW*�</{�x;��Ȏ�6��p'yh�*hW���8�%��2&EA�4�4�-=��K�*my^�/m��@/ۺo��4�z�%1���� �#�� ��)��X�[ZɶaS�M�@RNoLZ�k`e�����b�}䈥ڥ�p[�F�Xs�T�R7��oU)��T�t��H�&>�fna��|���ep��	��C��(�DH���pa��"�x�4pb-2�u����� �6�0�$�vd����
ǡ �R�� z�aT��a��H@���i��S0~@���P�$�9e��#�ʔ��knf��;�f�����QcVhU��#�k�Y3�2���R������V9}�H�*��>,5띈�D��J��R�"4�SDp���,�+z�rw�d3}��in�c���/�;l榄�n�|;?:�
�ӭ5��j�����_�[l��#a��`�Kq��.SiX�C����k�2�Zw�륣��#kC�{/���;��3ǌ��l��&N6���@���O�yf��+��+��3^�����b^���_�G+&�2�ȷ��1�D΋2#��v������`^��\</Tn�-�h��J���L�ə�9�pܣV�0R*����=�ٗ5���N^�$9%��0Tvx�M�5v7K���'��5oH��J�*���@!g���As�T��H-^�aa�o7дf���nm{�f���#8����Q,@���.>*��j؛7��۫\Oo�W��#X��#*�e�����2��D���L�,J�Q��j��h x���8&`B`���� K���`9#T����m�0�!��ؙ�i<�6vV�suI�(6Bmx�����Z� ڛ�aW͂�*|\Dnfٮ�S���k�[ �N�� Nr���97)�M:�#M�*�X �duCL��4�q@%f����[FmT��6���#�ݔGt�TS������E5�9�3�z.��B���(��̳��� $�[G�N͗�.�����W/z��M���؂�	!�a�6�G�U�sH��>9h)?��X|�u-z/�|�x5��t�)�6<��p8�U��y���3��5X���p��'�Do�"���e�F��j5�#���fE#���rb�B1�����8��Ag�~G�7�yB5�j0�xCˏ4L⟯��3���k��J��wP[�u_J;g���`k~l�Ov�xCAow}���ۡg�j�i�4��X�K]+奃uQ���_�l�W�ѬSQ��/���$��e��,�q����|��<5ά���8�.1ۊ��\<�Z�4$Q�/�
r�-���� -:�T����ދs�E��F��&	0�3�+\����Qt�X 7�R�X0��,��Kv�S힇j��rz�7rP�����(��V�f�%D$���O�)gX�k�	f�$�,+:�������Z���O��7D20����J�<Z��B"�@
�ɠz�kX,N��խzj�G����j=,)%j�b{C�z}�t�p	:T7K�
b owp�dC�<Z|��i�S�և��f��
���B�S'ڗء�Q��k��	 �`h(�w]v�^��a�ɺw֋yǡ�6gr�׊z���+j0 (��++�*��M�?�t�E���D���A�n^ν䑹Y8ֺ$�6
:ۦj���'^3w)�$��|�r3���c$E��ȍ��<3WԹk����:0���� �:VŐ��}{�B����`�Qw��ޘH��'d�"��Y�`W�駧N�bG�R�Ru���%�9ې�8Ǫ�X�F��2>�QY�Xx���r���rN������Յ�J�$�uʶ���fftA2�s[�/6/�����$z��i�5����GB#��BR#u~)k�����۝��[R�Gى0�<6����c�Z��.��,P�2(�?I5�����SYؑB�rRKn=�g����Y	���1)����!s��!������ B�)��r�I��&�<���^�`E����ڝ�mh�,���lʍk�rj0ڽy�����ů#�?Lr�u�[���'!���\Q��R�]��9@�s8���#�)eI��0>�[:pj�7T��!	f.���N��
���J��rg��g�0D�X��x��v�w��&]?� �Χ�E�y�~�Y��g6�>!|�81 ��̲>Z��]�<���]^ܴC_��O�m����&B.'�ԕі�\ܵ��
� }�:vahzd.\�9@������P?��ȡn�s���3����3u@$ْ�2�&����x����}ص���&+s��av;GEm��?!(1�e�5WLMo/kL�9NqXQ-�5������|��(���6R:"�Q>EJ:��'dQ��0�x����}-6U_�p�e��I��Uf�8O� p�S�:PS>�f'�@^\$��WR�zeg�i��nǾ�iL�^p&Up�L�P�*s�lֹ���k���m�T���e7��y`Հ j(�>��ōA���q74��,����~|`ͬ�z�(��@��+�UѤ&0�婟L�	�:�A�@ӧ��=[�Bd���mD��]��AQ��7��:G�F� ��OfC���壙Qr��/Y�E�g�����j��@`�f�*/�k����o?��8P]?��!uX�xW}\NL#ir��'���D����f���<hP�bc������C%������^1��[3���e�h��[H$_-b�a��7�A�e3 ����0L ��1��[C��5�ȯb��7��y� �Y���� �����̛Y�nJ���AW�`�z�3�\8���5�@���)gtFl����E�4rM}g�*I�Ѕ��(����pw�b�	�������E����\qtv�H8Ҹ �%Mr�������R*�a(~=��U�Y�ySߌ��!��������U�xwv�����=Ea�E@} @Q�G��;-�	g���`�b�$�ho����X<"��A%�yPs96�~zãY��5��C��
�0����T��h��� ��3']�!`���@X�f`�RZ��*t0Qaz0vp�M��G~x,и���K�e�a�6��D�1�D�L;>�O�>e975KT.�ß>d;����a ��ɤ� !�!<̚�;[��Wb��0�$z)��u�?��v�At��(»��Q͸�t����龏�<3����F�Xrm{���V�B��������4`�7d���0����4�-O_��ozˠnf�ͫ0�:��I6�l������e�(���%����^�|~���*�D���Э���c긿,�nόy[t�k7���l�PL)g��@����@�`�@�05����C�_P����C6�[�,��g�:����ܞ�Z���C8�2�]����Lz��[q<���<�@>ԧ|��]
Tk���
�v�@�8X	׈�*b;C��~�(��=��I�Ã��=cnt��9��e�%
�!�7�oԉ-�����/ʒА'����*}��<Fc��B���z���y�6�c���	�t�r��,�u���8elJ��2]"r���������Jʭ5��?��osc�*�tiA�	Z�!C���>Ze�����wP���8����Aq��{n�yŞl�yX����M�1vݳ���-.��wE�}֋XM=v5�ʢ�E��<8%�T�����|��-����RhK]k��I��J��x��]����Z��Cų�i6��i������\� N���.1eӨ!o��pWv�AT�梏��da9K���Y���*�x�j#}ܜ�+�1ֻ:�$-yg�nM#y��|��(pZם��rڼ#ׁٞ���Ӡ	�WK_�~+�}�IO?3�i�}j�MZOG��VR����?�� ���j�`�уĎ����(_҂\�fb���J#�iv���*�v���l,��E��=&���}���v�4��E��<���sf������n�$b�Pu�/	%D�p���8�g��=�N{�֗���LN�;��h�Ĝ$[����_�3P����qY�w�� ɿ𬾽��Ɯ]Oi�	� ��=�3{H״d9�?�GOB#��B&�ٚ��u�:QV�w�u�pz
?1'g
�5�Q�C��n47q�ۘ����C3�С[�(B���@R�Us��"G�K�^�4ʦ��:�ӱ�����p�О2�]3�׭�v��}�f��Q_j��A�SS�����5�A�dI���@� '��\�?_