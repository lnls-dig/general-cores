XlxV64EB    7a89    15d0h��s��w�f��O���A6�L�g�P�p����0H�IA�(j�l����-;/F�5[�ń�>
S�[�J�D
��-��$�4=N���F��)��K"c�� pPz���̗#�-~:bLc���z�M�Ίi�����'�d}��� ��=��zO�I+&.��/���N�@'Q/��$fe�/�fQB��e�ۋT�zh�O��T����qG�Y�8�H��g�nu�<�P՗�]al��yg��f9#��K~	$�������8@"d��B�2Ѐc���y���)8��T��/�P��-�.�ǳ�P�~��Y��s����0�@���� /���+���/.�O�(�i�F�Wd�ܬ	F��4f��N��_�b��F��Ni�dd�� �%�_���n�}x.�A������m$�����@CU�Lp��C���Hõ������q/���ʹ1Z�Y�Qw���q��6�L𛚗�8�'`�h��xANZ��pcܚ�)�p�+���)����2�n�F��NRxs�k��sac�X��kmO��V����T(m%�~��� ��񑱤u����u��T��ff�Xk\���xt���N���K6��z)��b=��]��65�Ln�97}+�`��7N�S��e���K��S+��!�8�R*@l��ЊQ�t[�C���;m���v����f~9�<�ą!�V���>��)D�����+��ؖt{ �雪>~ᛃ�P¹=�Ay����$�3z�p���3��B�AXU�u�JT�b#��/n��� ߌ@ʪzi�����Ǧ�/���
�j^)���G%c��� E�Z��t�L�M��g���4?\K�!�����߀ٿ��?)��,��&2�:�|��b���U�܊��$�Gp��䆥�I5#m����Y���ye���K����Z��i��K�{jõ�racn=G/��?=Gp����{M~��9��u�(>�ʍJw��^��-�p��:��Ǻ.�L�ЕX�&�����i�2�WxA	���{CA�.Ik���q&,��c�V��l W�[���h�<Tv�*�8�GZ����v� 3��(5���v�Y�p���6��^�5T�Iؚ�Lqn���2H1$w�p%����S����eO�D���{$�ƫ̲5T�0�����"���w���F�f1|<Hޔ�I;�O�Fs���G��՘�u+d�ּ	��׀Ü�����~���hD֊�1j�3+
NToQ��Uy'����0ZgH�&��%�/����hs+|�c`�G��
x䞋�����]��m=D���|uN��Aˌ"�|U@����H%CGDth���^��Q����I����K��̅2W�Ȯ_����p�Wa���p��)��~O��n��k�ntYYi^��'Ѵ�T\0o�{2�&0!���䆕P�PD��7���$����/�Սth�qo�^b֪��0��>�����ԛ-;Ⱒ�d�99,�rN���i�Ggz���v�9��w��Q�k��ټ� �.�t�,e��gҸ�P���k�a�l��>��4�,�H�ӌZ����`p>��;V[T|��|�L�+,)+5�e��z��s1_�^�1�<]�Y(/P�T�=�-���x��o��ބ�B�/�K�W�-X����#u��aU��}�E�G?P�O>���-"���`���� H�)�f(�*ۚBM�e{V1�Æ�>��!V����W�L���M�Q�Z�=)�³�)��3#l���>�/g�l�{�9H��|��B#Wu��/��ϱ����<?�q���̒�Ǐ�)���y-�8�6]�4q�(&$���������{�/d��_2|MFQD���$)�c	�Y�IL��.;���|#�`Z5�z���&���HAz�]����vK�2c�E�?@;��`)��J��cTB�2�<!���5�nZ���E@�I�����u%�8��-��w�!(���cg-|�b��9��}���>� �0FIW�N�s�\�IY_��}�
"��\�,F˓���$�{�C��t�>�y�6C�Ӑ�!���������Q�	�AWR�A^򌺅^���q���Ɏ|p� �E�U��lfH��SN;4���8�?dz�X��B����0-��>6�-�>;&)g�$s�x*B�f]�3���n�Ł>4}�.H���*3&���}����c�񙽅�z�?�3 ϙ�mw���ތ��ah/����@Xst檯�@���ρor��f�eO�;�o����W�,�a��������1ft��/��0���G�v<�	��wJ���}Y�]A9>?5�k�j��FSl�����<�������>G����m�T�Ĥ\���;��W��cDGc����[RИ)�����o0�;y[�/i4Z+G5�1�䒬v#Y���i�+�E�QT��ˉX<ߛ�DǢ��$�������@��'NVt�����G�jE�����f�k�hџ)��m�PGнp]��g�g�G�5�o#��Lw����E\of�J�?0w�Є��݃���A�p�8H�����=f��ĵ�8hDtS$�>���h�궧8�ǻW=�#��r<��
�V� ������J0�^w�r���gC��Q� ��W�G����T��u4=��N�0j�O�㪉o	��|˸�̓��u9J?0�xڙ2�Ў�B�|���[ZU� ��e3b"��sb	�Kr/��<$ *�k���'�2P�mJ���NG�{V�k�3�����?7ABE�����לS��
��J�y�����fY��*�K
8N�$�9�F����Y�ꙉ6�X�@���_�W��sZ{@�;�+T�B�r���٬�Ԗ�*Hh� �D�ٛG�wu���S:����"��I'�a�P���������,�n8��B�ʺ�MK0����d�Z?�Ҵ����:\P�fn��|x*�0���VaP۵�{�l�q�8�Ï��o�ò�WI��}$9)E��������=�&b��_����|�����q���t��"�^��b�-
����f��'��*[�tRE�Y��|�t;���7r0�^^�� ;!T�ٿ�'L�LL�jOIѶh�|䆊\>?�f;p��w4��QA�n�ҏ�L�r{2h�_��A����*��Ji��<��5ι��&��� zt��<AH/Q�l��p��9�4�?���D�gwwj�h gʑ�8�$���T�H��P�N��mJ�f��C�mss�����a��z��1]bKEm�1�剢����}���A]j�F��X�Y��k}v+^�|��CMݨs����>?{U�;)�>q���*Ο�sHK�;z��lG~q�|��3"�I�TLY���-�G��G�ԅ[��Mh%���B|CF������8�c�ʡ?*}�h��E���Vj���C�-[����BR�,4 -�����iv�D��N�q)�02X���Jn}��F��G�V��C�ye-����1���my��&�C��@=rxA�4#9��udv�����0;�W��?��)�[�޲ݍ�RЀ$�����������ru�;H<����]���	(�F�kNr���s��|�E��"�z9t,��-K��E��k�̒��Gґ_���.8#O����N��3� �~�$�Բ�2��έ�͉&����l��<����лu���~�}�[�Z{ƹF]~<_�6f�����;o�w�v�h?�l�(r��P�r�|�=|��z*)���2�L߿Zͨ�o0�dlUe��%;�o����~{�$	+?��V^3]&4��[zd�b�F=8N3����p�Gp��8ba������p:X^�'5��Tz�rYOE�z��yuM��gn��թ���<���%��� ޣ�2���[�zi��CS�$�]�g�n�z_�XVG���d�4k:��g�u�g�n����T�J|��
�P�FZuz "���d�6/��(v/�,�
��QS�E�+��W�ً��G��K�BV�U��f�ph#5'si���>�m-�E�Q�|����Pji�+q��0�ME[Q6��6?�1=�d��a��B�YM�aV�����Z�������麏�j�~�9E7�3���y���k�t��'y:�K9C���+1}Ow�0n~\r���K��|�<H�$�����	O�_󝽮�,��g<!��������/�ۡB�Dg�!6��k�'��`So.ˣ�Vq�A�rK����22&���q����I}��,�v�;��GD+t�H6�"y��D��?��J����j����2��L�>wj�w*�?>���k�zn����͞��X��D�0��B����D�&�OR����uB�2*��:��P�#�����7�e��td�U��S$*��xًZ�
rR����ȕz��W(If}"׈����I�RL)�,|c㴡��]/ �� ���S'����eR�c�o�'�I4S7���s��m��;�� 6��Q	`Z^0!��#��;H�=�Cx�6\l	ȹ�|�+�y�˭�D�.�U��&�ʢp2��Q���M��Ѵ^�R��$����;�����]�9x|����f̮-/�1��J
O�*\�kV�pr�G�K@/����ӂ��S������ٲ��K?�Ч�EQ�*�◆H�1�x~���KtY٘0������\�uLX�	ݖ�wO\ۇm�_��w����2ݰ<�I'M������m>җ��ý�@���+���:���\:��rh9h �cĆZ�6��&d��y �h!���D=޽l%:���*�^���S����������8$�%�xG���v�i�M�����1�'�Sؖv��B��	�P"��>� �Tf��&^F[)o�v��\z��F��BU��	��Ia;Tײ���؟�a�u䭍Ҫ7O!�p���*��QpO@t��^��_�]����:=�bby�By�F��C��D^�g#߸G?�h�=S�g�]���Z�ɟ��|����\)���U���ͣ�{�U�5�⮗�>'�A�Z�l��V �s�n��\3Ǭ[�
>x���.��}��lTp�zo�(tcU�V�!I�'1�(P�	�z��U(+1�_lS��~��Dw��^�{��z�֞?����r��^u�d�n��f�C��"N�qt�+n�:nf����}�3�0��g-#c���/@F�`������Ht���kGf�F�P�-��!�΅���8�nJC
(�m�3\3�A�Y�� J%K,��m��N2xKx�Sm'�?� ����eG*c�`8�?��i�4�J�9S�C���V5�%�,T�Q�K�t�Ŷ�OD��B�R�O�Z�#$q,z�H�2��6m�,�κ��E���4� v���J�F�p��x_��`���K��m�}���,���o��]C�X��Ir�������rb�H7����������ԩ�~�>�����S�T�m�8:��r�X����%��:
��s��M����8`�U?���`8�U�