XlxV64EB    25df     b00��*k`�ER��^�~xL�%7	��!Ӹ�8���M�@JTZ�C+x�G��n�)��7?���8!G*���0�9:HS�:Ly�8�_Fy�%Ml����礼N���^]��qs�� �v��Z"=,�ն^�k�BVײR�0�����\E��S����~�?���\:�	��H��4�^�侬	W�#��rcQu���{i�s���>���Ur�ݻ�f���6or63�9�T��I��Aλ����]^s�<0T퀌�ǆ��  H�QG����|���LG��(�/���IY��28�=D$1�a��
��H�/�t���⦤nBݦ��k��ܴ�A�mkMۡm�h�s�Wޣ}q����0aM��<z^�������g$���MF��������1]te�Ś����N�G/&{z��G0�l�ӆd���h���9�<�F����m7�u��5�fT�y����}�/w X�F�B�#_ح��0�jY*��G���A��s}��2t
�|Y��j�Q��f����V�r	�<,����ȗ'L !!�`�] ���+���Wfd�#^���_�n��N*�5�# ^?:]�k���i��R1"��;�/W� b�4֎�M���X�-"���	�������T-۔��L�s�.�~�-��2KZu�4��Iv�+�@{����o�?�3Ώ�*Dz	E�W;�d}���̹_ӲAqq/�z��Ts�f��Y���|��\m3"Cg|�1)��#T[���7J���	��/�5��^V
�b���LM��(�wʼ7�����Tae���c �2��u�<�b�VF�U̲�~�tA *���D�r5�a�P/��֫�n_ۓ���t8�3�h�[š���ț�k�ƛJ�6w��ZjM'�e�%(?�*��J	 /+����nbE����\F���h`"��h"7ev�'���D>�-���D�k��6�,���%�p����NW�X��h�`�^��zl� �>�P�f.3��n��49��� V�F�R��}"�4B�72S��:|�n{�����U⩙����X������P�4�Qu��ٔ�Q�o/�-���8`�r�"E�u�ܨ:o��E ��NU�`����O(+�0��.kN[���`�YTM��a1�MV�p�J�ҿƁ�_N����IH�N#�NJ�8��S��A�]�l����W�FI��\�NȘ6^�����!��n����%N�JCl�"����>��)Vw.8l| ����v<�}w��o]*^7���@��Dh0A�U���i�Ԧ<O �B?<�~��K�(���qv�ʪ$5��D'���׿r$MaL��n�	�>��*�Q�m��қiv3�ِ^���v�FN���d�/�B��8�ٱ��ޭ7.4:�(�D�
N�K�f�.a�Z��NW4�l�� �����O���2����ݣ$ka�3=y�QAA �\��(~^�-�	s��=V#����I�g;e�����;�ï�/Wp���x��U�g��9<�}K�"�N�K�$:��]O!�.�6�r����E�������W-�Je���{	`�x�hp�a���(�귥�t|� ��̤�?P���Ȥ�ݵ�`~����9�Q��Ol�Ry��dP�$=�j�@}Q�6cW��ºv�q���v�u�=׾����CsZN׾25LVV��J�h.�4�����\M����Iy�O�DY�H5l����(�~9���JNT��Ɂ�;@#����G=�Tai�τ6�Pܠ8��1p���gP����2�*�I�i*g���/�����U�d0��d�C���v�7�*�3،0\�hB���u�?Q}�e�8�M<�a,r�Nxjw�fIӘg��xS-�@���<o�&�H�U�5��=}�̜Gq�yi,����o<H�>ѣ�d�З��hf��a���m�^�!�twXKM�F����ځ�o��إ��3TzT�*�)��-ǜծK{��G�ߒs�E���Y@r�V���\��������s�TAG����s�n���9�d�������g��[pϏ�;yA�l��CЯ�����+�8�*g<�����׳��b�=�n��u5��0 G���G�W
�Om�
[�%v;���+�e/�@�'�Jʟ���5l�"�$�x�e�6;.���Z=6�0��Sh^,�&&!��%������Ū���jM��Yv�(l�}���t�]#"��Q$��kV�`�T�����8K�
V�����}��E�bYP<�#���[�N�����S~��'��*�0�g�'u��9Q+F�o{���q����13�}�3�K[-xg{�f^3e�s��/�4�H�3���*���N'��\&޾1�w]���L9��k����bˬ�r`�����p�R�]�փƯ�˒�H�๦
���,&E�?�~Ã���<%���{�9�ڃ���:骄Kn�KJٮ#ܠ�c�M_�tI�ʛ�����k�$۵|��`p��ߝ��h:�+�4�jǎ����Vȩ��=���iͥVt����I�b1&CE�(��)�˙Q�b����+����9�ܮ@��r/'������q�g��Ӧ�п;#���s5���>=���~��*�p��~Hnͪ/w����3�Å�^� ��l���	yT�;���������H��n�ō;�SZ�X4>  �ZXIӼa`[�F�!�w�ja=�">�L��輒
Ɠ��)h'��0�A���oZ[�~�q	��*���]�QSϟ�uc����iµOL��j�8lbo�