XlxV64EB    2580     b60�K=��j/�2��{���<2�a����GM����)���ûb��� �O7�Hs*��}����!��'.i��������׋̢�8���A�����^�����-��glj�-�Fd}7m��Aj
�B��{��x����r==����~X���c|������y��6��nR/�͂�쿽#���yF�V���Xv����	���n��I5��������L�l��ļ�M�����I<�!!H<��J���qW����܌Q)��[�č4~�,�k�������T2�T4�-�-Μ�t�9@����z���cX�x����yxE��`;��Ş�BU�¡��^��='_�0�6cz�6F�΢r�iG,p=�c���x�j4�)���SR�r��M�e\�b{o��&�Ͳ��K�4��a��@�j���X�TF<��ې�]G�\�7��������*R��f��XੳDU�zm�\�:���0�\�ճ�N����:em=]7U��b�����,\�8yK ��9��)ʤ�(R��ֿey�oc~%]�鉮{c��;�Ǉ�7�9����Id4�S�� ��9&�q	��� �ց�1E��\
�7k��r�=b��uD-���T�f����?�[�V��Hrgh@�F"k�^U���-i�f�͊���O����x�����f}0��A`f�ӟ�a���Z��V�\8�0m,CހO�V<�%�^�([\u��hR��أ����(%��L{��G��$��\��j7��W����7����%0�xGl��g���p'����KO�\,2<[�D�*��&�ki�5�:$��I�[��n��ػ���RU�' �%T_��?�Yn��������h��Pj���F*�][Sav��^���oT}T>.�<�v����;�w�hܴ�"F\�G�OZ��Fd��[�<�����5E�d^h>�5���T�~"+'�r7�HJCLtԢ�S+Ɋ��c<K|��m�JC>�o����4���'��E�	�!,G�4���k���ji,2��
7D�s�-���2
gN�^��Q�߄�}�E��� �W&���^e8Y;���r������!��yTN��5��ԣ2�@^���i.�;�U�j�a�Q�ey�^m���럾u
�����v!��F�Y�|�`����`b٥ߋ���̦�g��.+L;ǒ����{��e���O�D%��y8�VyQ��۾ RU}�oB����[�I!u.y�C�N!���Sѣa�bX΄�U5t~r߭�\q@塍�4@^�c�`�E/������Ѭ�ns$5�1���?~�Q�����o)��m���x#����V�Tq���%6&:g�����od�����qB94�T��>ۦ���y]�Ž�`�7��ebh��F�ӈ맹�6�n,������Yl�К{�RA������k8!����5���N��I]��&(�N�c�2}5(K6���1M����7�_���
y�*R_��1�q�&j͏�(��S�d�n��#k�m�����!�-��&_�)�Xg\�$�y��������R���k�:w�C�Tv�&�9�-���� ��v.��3���+��a���'k�"x�S�nVTMŁg~�5L�Vw�wE�3iw�9�DJ��'ܮ�x�2�i�oR�"�'�ji�>.۫8���ܛۍ��[_�h���~����:�H�<i��Ĝ۫݅WXW:���Y��뎸������9��zv?)1M:dW�}.�|�Q�Ü�T�!��`�|��"�I�To��-oٖ67�ڍ+dw}�h�|d%���k	�a��-��>��JPn'ǾB��_'�-��ƨu��ڂ! #l���9>��z=� ��o��^��a�&q�"gԜ��qH\����!&+��D(��6w����VoX�jD����9Ұ9��j#�
��-�U���7�W�(O�Xz�oO(�G�@�����l�?�n�>V���	4����گo���6J!/G7�ƃ��S��@�x��
�;Fg7:4L����c�(���;�0�T�{2�)�]Af��`�]�b_����$�DxG���6�R���NT%n�K񁿑^���"�h��D��B��Z�Dr���=�J���GÌs*�̰�
Fo3J�y
)�WR��Cs��P�">�y
VqRM��ʴH�5Ԅo2l��z߄�YI������í�'�x�qG�"7�E���d�r���E��i!�����	D% 譭B�70}P9T��(7�+��A�@��B�$M�wB���-2�g�kE���
[�bT��W����
<B7�C�k�w�2U�ၓ����>WkZ7��|Cq^d*PĆQWY�I�#�D1����Lx���v�+6���42>%���@�^Irl�?1�UX�R�",-�� [�%N�����S���ywG~�`�	�Q�U�pp�mcoI��g�%��wH��[�ƾJ?!���v� ������ꐊ޶w�R�I)�k�ݗ��d�9ƶ��dK��'�`/6"9�ʫ���GS.��ڃb*��`�Xs��@�d�(�mli��
�����Ut�}p\�Gj&%Nbm�f4ƞ�+l������KC��8�a�j'��Q0�v��@0uqFF�p��+���+R*� '�|�7`7$h��j�P������*�=����	&�l$�'�ɹJ�^s�:�V�Ƴ�#��"��nDQ})QZ�}Yh�6�)I�������ݦ�.*�qa�����Go/�Uvɋsq��w�ly�8t����\��Xѿf�P�W�öFۧ`�MeP۠��;��	E.*�/�*�t��nY>�UT��ީJ��C�O��M�a/��3�wE��P����eJ��s��'��*