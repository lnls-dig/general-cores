XlxV64EB    df84    1e70���zm-�W�y�ӈ��������s��c����_j�/�Y�+c��c]ѱAwf�xh�	�=���Y�msb?�lO�B�+��FӴ��'jM��y;��K7jn:�,85Vc��.�AX�-^d�Z�Em����+Mʣ�X�������uq#��e�^�=3��#�ޭ�� �#��$�\�2;V�	X�|����.j�:����wZ�Ψ�!��L薷�~6Q`wLIk�T�$T9�(a���Y���j�J^�|�b�`~,���ɐ�*� �=�z�����5Tٟk�:yߺ�H����RC������ ��:^fH��	��5���B��a�+�Q���g������f��	j�Q
���K�=HZgF��wU��F���U�q��r�2m}@�(R7�	Ӌ�|��ns�.�E�X��_�zi>��&�y֎gP�تg�=?��Po��?���z�!�����{YF�D݁��ԘU���� ��'J� ⌘�g��L��X ��~��Lw���O����m���~;�֝lN��f4��ݗ	ŮL-���#J�lhp��g(�)���A�*U�ᮩP6u)��S>�C?3�ہ��\8-�(��"�Kyj��J��,?E�Rh^�$�����l��P����h�����F�Q ���x+�1��w���)�3�d�J�0��A��
�b�*�	R�]��Bʞ��դ��3
>�P� '8��F:<*[�����ЂVH���i�,�0�8�X>w )̒M�Z@[��k�]u6f�u,�eڣ��}�Q ��3���>�IS�3��9�6�0�� ��BZ��oa�x:k\�l6!\��� dD1R�1�?֊k�0��|S�fm�/?4s�-��c�uQ�D���B�L���)BӸ5lR�)z�ER*���4�\tη�b��J��sS�Nhm�q��\Q+�-s)K�
�[k�����ӥ��$1���������E�������&$:� �:�L��c*$	��M�ҺPEwG������M�)�oE9ЬK*4�4pA}XO{�9<z'��E�{Gyn�E�G���.�vS��G/��"_qYL��X��g�xȠۑ-{\rSr�u5��.����7�vu{�s����L�T�;�(��W/o�'RrO���q�k�F�Mo�Ye#�՛�,�U`##�Q��R	�EyMVSm	�QY������1-3Oe�^К,9L��!O��w�[�P�P��w�!U��4H��݂;z~���C�Â��@V��̗}Q7�B�:a�6����0�av��\Ó�PG��u�'�1���`mL�9�A-��NZR}����3�Z�!SO��d��5��W�4���\�ȩ%O4�+��>���+��8�<���ֳ)�F��d��^a�`�&����t�-���Q���V�v~2�W����מ#����	j���kQU;��]Wy�؀�6�aj��g�}x�z�i�_$J_T�+}��������Om1�&EDF�n5���K�1*&"&�C+�n��<e�#�7�
������LNI�ڛ���Ԯ�}��op��VR���%SC�2�,��v',�G-Ȧ��G[��R�3I3pk+��
��"��b9�.xz2o��Ym~����t��P] �鍪�5���ǒkNh��y��0�_����y�6𾸖��}��~5Ӧ��|g�\јf�@a!5�J�x�'��[�aU�!��Ô�j$[��p[�@�H��v�87c���o�{?V�"�Q6
]/m�w{^@� ^JQ��u���"��E�y�^�p��_H@��b&����18�I0���G�KGj�����¸V���9\�m�&���*�D3��Hɗ���_��T�G���?QJ��e#K���[�7��%O�%M����/\�/�/Ԙ�a|���f�e�RV&k�"�摺�*c�� ��JK�µ����$3�1��A0�sEC�e{~�;��PpK�}��m��H"�F>���ONW\l�s� 7��Z�RA�.|E�1yͿ� #Ʋ����b�g��*������D{�!����� ȑT�g��=����*�zA�t��d�z��Sj�a����"�k�+経�)l@�+�f����6�R�OKV0�^F�]�\�u��{.	4��wb}�	0'�����C��~7��~�{���b�kZ�>�O��ɵ'��2OE'�AA$'k�Q�`���VĳR��Ja�t�P�'����ۀD&�LP~��	����Y��R���u,5p��s�F�P_ʿ��Uۭ�܍�ز �4]�U�vo�����L�Ȭ�'N��w�3�\���u�� �:Q�6T���[8�����T�vB�&�����&�T3��O����U�}�60��S��/w}��Mg�H~��X�/��sls��c�G�Fv� �!m��B�V��d�i�5j��\��q����N���B�zi�]�.1I*#�E��h���"<����ң��>�>��g��hȔ7�(61n�x�@I�9��Rh9��	ʣ_3*R�b{mb��h fh��}?Q�!��#S_��:�FBm{V�_��+�U�Zm?�14�ǣ�T/��p� W����1����βB��N'��Y�	Bp��Hi��+WU����}>͆J^8B�n��/����g�V�8J���^܉�K�m���[,�Ti.Y�z�
5�]�y�ػ�}�[�#�+�O[=q��Z=���I���ew^nlG�٪���F�
�Є��Tci�5����vz�r^���vA3��=�����>'Rhl^�j���.�	6t���YC_"��\���A�R��oXd�/�3ϔI�9�T��b�B��!��8'��F�㟘�����)�~�Gj��'}1f�1L8���u��1>�s����ԡ�I7y���(�O��|��>n��f�_�_ V�����EV�TE�k�a`��5r���.@�B��<����q��Y����~���о;�ԩ;:�?��K��Ϋ�M���G3ϳ]��_�`3g��)�u�I����}�i����7�sI�/�Y�D���J�ƞp��d?e(� Yn@(	n�M�(õ�N}wX�hB&���C�u��q�d�2���zQY������[��b�l�&��(Pz����i1Xf���Mkd�hE�8���Zo��1omt���x�-nqv��������5�y����~�V��/�1S0�+ ���z�xZ�y�5m:
�����BH�MvE���[i2ذ7��@dS�%^�z�g����7��g̈�`xQ���������4��$���4���:������ƭ��2���W<h�'��P �֕r{����ڋ���0�oF���0Dʒ����Q+�P��{֟H&prͪ:��L^���������P�5W�%�h�ж���aCw#i�*�9�C2�8�@Z�6N\[8{t��1�N,9�H��<�T�cQD�����HS�!��s0���1��-���쀲�eN�v���K�Ԛ�Ie���'�����O���A��ڀ������;���œ3׌\5����.�c7E�x�a?�ѳ$	��j;buL�l���|Ε���,H�}�R0���_���+X����ɯ�E)|���{����m/��O�z��Ψ�,R
Wn�.��Rd��v����4��}黻FQ��8�8[�'n!j3mI����^!֡���`t!G3��̩���t?�p�B �c�Hj_hN�Q�a�A�/!�
�R�Xb�L'wNg�Y��DG6����� ��R���mE'���J�e����.���՞yK�e��{a�7�t�5{mO�o3-��0��	u�8��pu��9-��i"�"Ƌ�x����N���?�K��"ƜQ�s$����`�;1S�������B��
��x%Sm���c+޴��(��7�N��D��.��'�%���������s45���	?�s�fJ�@]��e�
b+�h�V����U9^,U�鲢�w<c��y��:��k(��n��*x���u� ���;���,�f��*�95L�kUܩG*��v�+���1\X�ܳ�����^F��=��;gk~�GH�R�y�B�vƅ��I;�M2��b��;F�2�KF[�<N{]�/Yz���*D&���QT����s>ǝ:���O#6f]P�v�,����hBx'����d�i���5�M֪³a���<�}V�I�BVv��)������Q��!PW��ڈM�a/
f�k�@�h�V�y-�$��[.�]Q�1����	�V��H�,F��� w|��� ^�'
��(.$0���;NG�򁻛������X?�-��L�i��'��vىe�z��n��?���ѴU+��>3��QCi��:����2� (+��x*�/Z�������c�?S�*dy���//��?SH�@=�C}����խ|$�N�����3��A�l�4��ߜ�rk��on��!�t�N�_>�F���}(�'N��E�l�
����t ��*�hO�S7�YtY�0�|���	R���K��68p���}u�b],��������=���~�w����]�=6BQW��W��Q�Laכw��F6B���Yf�d���P=}S�a״�#4���'�o&�w2Ǧd$�1ǘ  ^��̬)���Tm�D���wޑ����3gh}���3|�8�-�i�)&��@V����u��Ȗ�R� #SD��
�!W�,�ZV�/D>����i�q���?�V�ݛ��Bx8�$�eJA+CK��Mo)�+��	��e�����Or��C�}|g�㨷�\K5���	�UC�����p���BFd?>�� �[�`�4X���)�I�H���]�y;�U�
�y8V�����[�3Lf��c��<��F�5Y��r��N'�;��IY����d��Ft?wuiTx���aQ�@P�@����>r ݾy����lJ�	HP��2Q�춊�<gpk��S�8���~X=���%J�-x�ű�h�W�㘞^i򺇠il��=X�s�(!�o`�;��"9a	���g��4�����I�{�j`^?���4��^Y9���`�:��J�l�U��}o��ta�7��-C�����H����F�,�ұ���;)������Ϋ���մ�^�te����;V�3|O��.��r�6��v�'��\�ߦ�~0�F�>Wڈ���3J����Åb���Q	a,55����oF����^Opuj�{8�����"����n.�mW�y�>!�Ku�"E�%��&��4n���b�%T%��=r'w'���f����p4\�9 a8lv��vL,p�|�[�-�zZ�ƄD64�b�m�n\W�d�G$�&�u��b!|M��\���U��VP��:EVM���1��D�6�JcО'ؿ$��,�_�x�/k��z>[�>�B��֊�����ȴ�.�l�dd��bwtu����%:r<�2Y-�Q��{��T2���I�(�d�dw͹%F����u�����F�����οXw���J��oz�8�g���ל�ų!M�-ݼiH][­.`/o�D'!7�,�1`��댑G k�Y� 	��>0��.%�-���$N��	�U~*56C<7���f��l8��?�R��_T���	�8٪�1f�iz� ��������9�Lo�@ G��|�HZ\�M��:}o1�0b��Ȑ�A�a~{]Ӥ[a}�_f�[4�:1�1�O^t��}�V=h>�o閌��uT���|�cf�����7%j����
��IyM7�D8S衹�ȇ_h(�PUG�g�'5;6�X5/?`N�G���� �X���ЛG�����|WY���g{u��oy�p V�� �5�nfv�zC���#E�GM�zJ��?\�zm~I��i����;��3=>(-l������+㻣��W��f���f��Z�!�9��谉Ea��2���a���K���Pl���3ܒKL3��h�O�l(�	�h�
��J� ��e�秵�w��Ϻ��Nk���&&t+�膅ʷ�����n�TE[�Zt�n �Ż��������%Ņ�1���){��j��OU!�/��vl+N��ZJ�Jǥ\*;��	���}�<)��pͻ;]X�a���&h�F�<�`>|7��G�/r&��</е� '�^��j�@�E�?�B���R)�h���)o�?��I[n�?�����'�ۀ"��,(r/�%��u�)���)[7��u΂��`@p��AT�X���t���
C�(FՄLR�ZH����}=����X�Jx�Q8IDbQj9�Li�pKa���@�y�D��Iz,oiF�~�ma�3��-P/�I򢀇4[�!�0N �	�s���	z>dL���6��=�u����o6�F��ϩg1j��Y���͠R[Z���4�ە��V!(��C2����ܽ�5��h/�) ��!Ҽyj� ��3 �ܵqdh?�Ӥ�LjYX7Om2�w1�!$�E�h����)�`+]����:�d����Wze[~�w�kE����/�t8�:D�����=�j/h�6�d�
��
�l�������}l�m��Wqw�ҁ�"�t�_各�t�����!��x�&T#Ԛ�K=3]pȥ͇#�ǰ0Q�KC�ȁ��0�+*d>	)��>����.T�q��w�������v�����5�x�잋�!�wQdԹٔ<��`��v����o[������K �z}�ު��%*v�[Z��⒢����Ol�wG��R���Axޔ�ߤΛ�Y=S]I~z�����rollĕ=b#����L����旐0^}��$	j��}i���bL�����3aW� �9D3��]2�7����',�!A�ڃ'8h5_�K��5=�{T
�����b_?��(���&G�x"ק��������Y���A��$�'�����p�n���{�v}�M�D��`oB�o��>!����J�����Ϫ�����v�T����XJ][+����M�~�m�'�Nr�^���~I��'!9��s�]���y-��>�n�y��z�!D4�|cNz�b[vˤ��4xC�1���ÝA֧���EǸ#����	Y�����%���U��`Gh�"q�5z�pEEe`i�g��Wk]��N�H�~R�p��X`� Dq�!�u��"H	���;�B��<	19Wtժ�XQ�=�y`f�
�DgP�Tm�ק��F@�v2G	�˓��_^��;�_G����m���<I�������Ǭ����+�{�/j�''�&�����px�r��"'z�����~���z�YP�^�2>��n�ȘT#�k��D��}��{Lb��� ��L�Z��Y�~L�C�	J�<Ac�	�4����t��	o��å����EJC�/0��Zr�"��j�#x�nT��x�c ���v��oT�Zt*K��v��^�p/>u`��w��h��B�g��L#�K�M<k������}�z���u�2?��Y��
3d�Fm�x�q%���o@�'�Va�_.aPK\ ��������X-��oЛ4�����ߨ�s 3��ɹ���sh��>�"��go��-\m]Ht|Z 8�P�>�p���	?s 	b���؆�`�3�5�;�ܔC�R)����;��ܞ�n7�w;���4�8��&�'���3��m�$����1����W���أ[�2Sz6.�^���]��㽭^