XlxV64EB    1fc6     9b0o����x��nf�)4�o�br�+�:��D9��qV�n��_Z�97B����6�b����l�-f���W��ժs"�oA��5�{�l
�`J�u_�y�LHz;A؆S����Ve��۟=�(�D�=qm��h@%�
/�^���4��h�{E/{�-����R���I�x-�Ƿ��U_.���%LӮ�\��\��%P��v���:A@"��nc:��:_�}���hc����4�Y&�H�9�(��6hKNXb�T�W����G�aQ�Jr��n�xF!���L����dn�L���,������%<�qGoP�x^ �^��K�/�lI�D���~v
���l��3](3�\�X@��A��+]~վ?ьN�W������V���q�����v�x;�'����P���K�3H�׶c̮��֊��.�סc�te\��2�?�G�������X'�>⚸����� ^(fD$��<f48u�g���=Aivm��'�ɸ>^]�TA�����̕�V������$X����)�&#��Z�P�T�,@K:e~HW �x�YĶ�;���4jH�k�h���k�&2�8,����[�m��}
aF�1�w��D����߰������j�W�}	yg�ᙏ�`wQ�|�єN�`�+���U��v� ��2:m	�|W��C� "j�T?2���^�k��	��T�C6���$b���/�$n�����,K�Qe66�x���y�ϧ�l�)�3���2������ޙ����#&�?c(�l�-I&,��G�>�<N���i��r�W~q�c��͟�p;�����:�];����Z���Y4$�"����#D_{3?�X,�3\?�9q�,r|6%�E����[o����N���e�Gx�W^4OG~h&@hv�o���H�(
�jOu�;�%Ǫ��ixr5�!mb;]��}4[/�%�D-��E�6�]���.Ҝt�n]j�)�a�h,�ۚ]�+�A��A��*\�`O�w#�yG���$��z�/��<6 �2��%
-a��T/�쿢��Ehj�7� ;*��WH09�l���=�~�^ڛ9q}�m f?>�lь²��C��g%V
�ި���b��Krr�D���>�2Q��C`����u��0W�nsk�4ZhO��}{8*��U'`������P��C�>�k�	>V�E&�w�y'�N�����cr��}�X���۸������ZjK�Y���6<��NԮ���O^�$m,�˳����nG�/�Z�ثc�6�t��fi���O<9�ѣIuB� {\�ߣ|I{?2��z��S	[��.-e����)���\�sv�̦,������kY�������	1�t�z�`����rZH�����]�&ŝ�<ݺ:���O�k�e��W���,�J�<��oQ?т9���{ |{�}p��?#�>�i=���SJ��A%w���d��_\�p�3���:6L�l9��UH!�/չ��l���SmP�(����etU�y(��"�i5�,8�U�Z�[��Z��yY)���L0tb�=�m�m���Ƚ��R��x�K�|+�r��+��#n�lɂ_�O��n��nQ���0ȯ�|��r����1�DJ����?�JQl|N������"[W� =3t2��s��k����Dn�&C`)'���l"��,�C��3k�+4�DG�}�Iη�>�'D�Y�wQ�xx^.��>�I�ψ�ș >����m�0HGQ�y�O�yw���߱�N�G[��6�,�`�Z'�H6�	箩;6��X���wP�iB5Lt1��/�ON�c�ߺ1�2�ի����2�J��b�
�9�V3��<x�kE�y�qv<0�*Rgu�a|o��}k��Og�צ�~wJx����rM$;K�6�0����I8C������A����f��U�v$ *͛{�j���Y��!]��)�j����{
K��t����2CZ�u����"/@���.��7��ӄ߶*\�~
�PZN.�� j�E�eojnm��Ç.�jh=o��e�!�Ta�.�vס�V��f�̮�4�
�/��۴�\I�a'��)j��m��3�T�cx�UR�O�	���#A8����>USj��c�J��|lܒ�7pc�o�1[X�l4�28��Q(H�T�ɠ�z�DU��.F\���7�+�8�����io��z�_e��v�F��nY}#2��~.����dղ]��Ǡ�ok�1
԰|��ܲ���Z���'-��=g3��*A�,U��MD���_q��:(  �7�sx���~��#���E��"^��2z��ۨ��I>��d_q�e#�����g�'�'�_L\g�^O�e�-���Aa��v�`��..|.��덆���[��k_;^�ۮ�F