XlxV64EB    fa00    2500�����h2�Rn)3o�{�{�w7����b��t�%�t��?�Ѡ~��:'��v,���|q�~��z��w�H��/�t�V��z�Ӥ|P�c�h����ڴԐ�>���f|_�W��O&Ֆ��W4ڦ$w�[�����o�pF��ܶ'$7Wm]��e�k?4�G)5%Sj�:���od��hm����9��^��ח^�>+�u�_�qJ��"�cfDh|����q�(b*q�o��懸g�=Ka�
"��z����j�}�_����1p�������𸫌���~�z$��L˵ދ�8��Y����
1D��g�I{a~q�r��h��A7�´l<�eXB�=��I�F��`���)��F.\��p�t_���[ �M���Љ�F2����&C�pBS���܎��^� �����
T=�93��?e��0��S�E{-?S9j�6�l�/F^p�(�+�<^�6��:4�/bg4(�ݳ����ДM#�pmQl��Oz���79C�#?��[9V�d2��|R�u����&�?���ס��)I���� �EE�RIA�J���<�wp�u�����*�D�2!�M٢�{-dw�̨��_�aF�e� �*�_�[&�&��(N�^�T*�:�`�����mK�O���9�#Uf�踓,���2�-�)z��$O���%��e-r�,d��tj�����(͖����&���Ef�����ͩ;�*��5����E/��x�TQ��������CN���9�2z����l#�R]����J�_��lP������s:��/X�{��_�k�;��qk�n�,$0�^����̰SR}�0�-�i�����ig|��ǏTs�����
q��<��Rng	7wQ��#d<!���PG�f�����@]�Vut���Q�Dۙ�q�7�̐��v1Ti��OyF�/:�~���4�0a��?��|L�F�I��y^��Yн��2h�'8�R\��%Ǟ?��֖m����6+���ҝ�����Hi�eP|�c��qe�����:�O�������
������/�.�'�����֌���ԫ`4=��͏?�q�p`e#���|r�C��<T�9�a{�(��I�*��8�*ڱ2(��%�Դ��0*���sp��$�Dy����M�tdq[a�	�
 iƝß�"-;��pFߒI7Y6F]S�k�Mc��j�\Q����j/l^�ϻ���� Z����� �}���io�/��˴r�?h,I�>-�?o&���a���jՂ���:��.3�XN�������u����M�WtlU�ֺ���w�����L<��.Ӿ�c�Nސ����BXV$�m�OW/�����eğB�|O-�,w��|��?9���c>�h`�a��x9�W�x٠�S?46`;��q��S�W�D���8��}7�R�~k�ez�>�\M����+&��h��1�)��)t����������J�Z�V��T��#��j)b�ɋ>�!�J���r���1 ���o��ChfY[_�c;��+y�LP���$�ڬXe~BF�;�Cv�b�@�}T3�w��/g��<c�4Z�L�Í��;āc;��t�6\͕�ޠ�L�z�OIF,�14��0�������8�ˍ�z��¥c����e}U>9!����?Ц
[zd�A�w���VB���d��l��]wK�����d�|2�a��H'2�/�+霹0�Y�<���QRAE�?��j��	�#?���nz�m�m����V�%z�L&�yГ�֦<�r
F�ث�v�i����F'N�V������V�.��]��=��˛�u�_�ǆ��.�KQ	5����a3�^�>�R��r?q��ZvC����"�
v2�;E��@�hg�=��r�U�A�>�B��!S����V���� �uY�{H�x@�c���}J�oϷ{��u�J����G����Wq�!����Q�D�[����x��:��*00KWR�[���m|?6�T>iF1n�gt.��<�k��w��TB��3��[2n3�E����*UiY�K]����:���;
!�6����z��l�����0����W��AD	*+�{�:���%�l��q�CG���,z�������ı�3Z�> ������v���f�����1@ ���O5�ʿY��u��س|�{�&U2"���8�5�M�0�-s&���U�:�ڰbbT-5f���Ap�Ŏ�_�9`>�]j�v/��P�hХ���BDv1^CG�A�����M���o}(w�5�w "r�0���?��5�����Y�����`ؼ�	�
j��Ao���g�!�	HyJ�ČSe)w?�̇a��QØ��=�2�|VI�>��!�'-�u>��hQm��?��WYUh��:eEһ�C�&�����Z][s��ͥZC��F@��H;�����nɵ*�+0R0�5r�m�i���ǡXFNz�O�-�&NF?냜��"il�+�������oe�%�B^�����'`�l����'C
m�\h�.jC	�=�ŤUń�����-�c������� jtj\.�����@.>�<]9P�a��)�>TЈ�mp��N���!�a�:7R\��4�FTakV^���h�e������	�w10�$�$�BX��	�K[(��%?��g����~e8�]�+T�"e�'L;�}w��x��C��vQj�o��A<�&-��4b=�w����a
¹Y����Q���2^�Sts��p��n��p�,�m�z����Brz�֫*���I��^k��Gk��j.���A���t���� m��Y���2��:쓳,���F��:��f#~ap��a	(E�?3!�Dl֩!쩰J�M��a(�>����=��jnȈ3g��	�:D.����T6I�5,��9���x��PH��`�a3vC�f���(�/�<cN�����3ɤ��P���K�s��Vv��X�(�2���-(��T"�Q�L���=\�Oﵧfc΂pt�ϴ�:7NB�{���!�X:�v��Y�'R��e�l5���$�O�x+J��L��+���	�`���Ysg��k�/18����+['P�%$����N��5���߫���QMY7*�� �QY�{^y��������'Iҳ4��r��X��</�mġCd��8��AXIh��d��5:[ zP	=�϶�X��Jr�U��}�R�?�4�ݦ�@���л�+ G����?��1�ro��X ��q�NQ�F�+�̀���[t����K("�Ǧ&v�Ë��X��k���0��	n:�G�C��w.��s>{+��ۑ>�*c�L�O�<��/�M�Ɔ�l�A��O:.�T�p]OV}��\�뉬w�려�@�D	�����)J~�;�=:<j8�Q���DЕ���u����R������KVH�O�f�˄�ll��:��\��'챏��:Aɦ�-I@���z�^Q{K3ꂺ���q/�-�eLɦ�PޣY�,U��{W������b�������˹���*��Kο�U�G�_0���Q/ɑ�[�w��X�jE���"���L��7����}RS>GM���ݏ��xIm�F���m��Ո�c���z��+G6
dg�94�-����	�1b4��Z��t�+��
���O�� 0��]�;�����?N��K��%���[��ǉ���wv��β���k��ǁ[�0���|���yU�N(9���B#�����#\kq麨�N�e�K;�` ��z��/����w�x{����Z�M=�z�������p�N��Q<E�S>K�C<���"�BqY ���-��ݹ�~�A2�J�b���f	~���aA� �C�ρ��*ضG*Ofw<(�k2�y��u'-��u�v��"�pB��j+p��܈��۽ܢ-6��+j�w�����>H7�e[���W�82 �1�n�"��0�C�ڏ�-c��L��$d9���ד�>�w���6�W������-��V  ���_��}�Iu�kzg��&-Ds�+���Wr׬���@��@]].=��h�k�(��JZ@�_ȗ�P�_\Bdj�1ǎž�g!���=�X����7� 8�,ù��4\;�����A���� �Wt��Qj�h�菾nqTi�������VkY�p[xm^ǖ1�[O�����+�a�����:������4��&���(R��L����v��{(*ŗ͌�\e8'����XP�C�*[ď�FX�-��&��U�2-#�MrY@��Vq�.�٬�M���/O�͆�7p;?|3-��ߤ��%�(���>�W��nE�T���1��Q�L8�cj^?�AQ�xfJ�f>nK.�1���R�_J�����~����a}@�t�Y �qi3u2b�_9���=�әN�����I�t��Ǳ�3A�Ӓ�C��F���I�i.i�>d�v�ןobk��|>�V3�ZVSu��L�4���`'�����<ǋ�m�%1jV��u��eD��F�>U�3����q�bR;����li@y ���j9+��lIG�t�
���)���)v&�ˌ�]�����k�K��C-P2_L-�U.AB��i1��D�YqjX���ߙ_)�`�VP�(N��h����0ɽ3��h�81��.(����t�A�x�\���4��l�z��aT�ۗKؑRF��"����@w/^�tLM����J��of�32oM���\E%8c�F�`3����k^��D�܏�HE���k���R��J#�/>M�,t���P���.�L�B���k���A+"Z�N�j�z*\�]Z�{-�|����*�pO��9F_���(fP���>�n*�*���<�s? �"�U��/��E;��z�Ґ�!�I��C�g���%��Ӱ7���L���*�rX��Ǽ��'���Zk9�2h�a�H"y��y�����i�h>z�H�^G��p��ś��i :�Ƅ�
;a�%n�yD�ڤ�ޘ/�n����*�C�8[X°'Up�6����/�� ������&��''��8s�2N�z�&��a8�� ������!\�Aju`����*�0|�F��D��D���߹�Kd^D�L��ˢ+c�壷��&��F�uAL����[߽C�v�&Dq�
/W�df�PR��y�Y�En�.������| �J;C_W����:��7���`�#��4�D��w<UT+��IS��*����.���x��U%�>,�Vwr�z�;/��Bp��m�T7	��d&�Q�rquL�ѿ��?��)5)C�y���HqCM$@y3�*8���/$|�y
�"�_���v.��ǵM���I�:~�s�ケAߙI�!���R�Ϫ�m��6ȯ���*]�r����%ص_��X+ e�zZ�?m�N����/���
~����ܭ�ӑۻ&�¦^�A��g�X��S�1�`.y�1"�1 �k����Y��vI�i����=�땱�7�0ί��v��@虫�\�MϨ��^��;�6�0�߱�	и�Iv���k;�S�������W�=��ō���u'O
'䴵��E�r��1��g�y�M��u�7GB���on�?�~���^�2(GO"�y��
��<}�:+�	���a$��B�Z�����f����]!0%���%��V���R��l5;I"@�*��y�� _�R���#���|ŭ�v�U�<����r���~_��֮6��)��˟
p�>�A�
�i-*C�� �R--�Ct��+;�ǃ�)�GN�l4c�aq��ve'(i)ǕΛ$k�q!sVޣq����7P)HT��@U0�,չ������+rX�5%�N�t�f�ʼ��yH�l ��p"Hࢇ�Sl�Z��nr�)ޱ��f��n�����|�������K��g��<BQ�'�R�zL����ᜊ�o��W�l�>��&��$�5J�n�뻙:w�n��t7O�y��Vd��n��2vO�0��kp�&�F`�}�uo�IY��>��G 8���@���P��d�����j�\~�M�U_���]`�Ѳ�j#pŚJE��!f]z�	��Sۮ�P�g��[���|DR2� �i�����6��A�W���o"���i��[�P�X�(\d�/LaH<��}:��q��$Y�2��&~��f�b���"K��3�CT�ͳ-Ģ���T�Te�L��36�UY���tY����n�������:B3���寤c�n7!��R8��ez�����?>���#�$8�^p�z��7=�����Of��-�U[΍��0N���U��bMXBQ8>U/���/y��ऐv�Q,�L���MrbS�`ih�*��Ӣ�������8�������A���WՏy���sL��$�)]��e�a{*#�!���Vk�z��J���y"�?Q�/^����@1H^y�<Kc&��P�\��d�z�$N\A�c�L s��_���5�B���2��&��ϧ���G�脙4��R�E�c��*��FhD��t��JE3�
�{`���r\��'�~���K�tx;�l(r5�q�7!��f�u(�̢��R���P/Ï�� �v:����z�}77���$�e��ʉ��>�_�E�$u$�-�f����f���g'g����v��eDxy��k������,�Ӓ�7؇��q�9�q꣆�\�`�+
��D��1A
������Ӌ'
�bpH~	��vݥ8-�q���\��l+�z`K�@����2g�_!:+S��v7��GZ�f�䳌q�c��80��Nu;O�Wl�v��vd�������*�Q�GV��"�?I���P��������}a�^൥,�.����ʢ���is95!�.�L�v�5����h�.�u����J��JR�i�22f�h�O���Q�	W>�]Q�q����]�q��lHK*A�%w��۠3=CI;R���[�K"�q����)y�"�I�q��@��3g���Y'�Ghl��
��E�~�ɇ��2r 7?Ip� ��.ݴ�x^l��y�����{���c�����FL����ϾҫQ������XFT��{\ C�M�U#�,����f��F�Dc����d�AM0e4����^e����r5?�'���A�G`n$�N'k�ʋ���S|�1��z *�Y�`�_�u��[k�
 M��KD͝�����[�Oz:h-�iQd��)U+�� �YNx��N���� ����4T3�fS0g1�i��c��7_ClκE5Z�Ok�"��q|]M��8 a^�E�xp䯧7�ܨ�eꜝ�F��-�;��
�5�c�
�����C^)I�����J���m ��Iͮ�!�O�J��{���:-m��Ro����>ݙ_�7�R~��s���\ФJy�R��9]��������-G�e��8��<SMp��2� eq���eH���M<:��4�����|�K��*M�*������F+�c��*�so��3�z�s������\������Q����rߔ��`,��+
Cҝ�a,'�]y/�)B�ȰA\�U������OǦ���b�OWMXw� �7"���K�@�=2n�
����t=�g���O�B�ώ�1��#��wQ2��j=����g\�]uA4�����y�gR��'��#�O$;��>���� �(��4��q~x��;��:h�M}��F?������� ��&b!� ���lU����& 2O_�X�q�yEPT;&��*���"�������_3�S�<CKI��,"�Z%6uCЁ��������˩܎k�K��2�����%�+�`�{�pl0�ЗzD�f�.���];�{!R���ERN6*��Bx��t9`�O|�Ȇ)����^���3�a�&:l�s������9�CvG��<��o��E�**y�Q�2��Uv���kt�!28!�Q�h��VFɼ)cf=�^��eQA:��"�`���1Jc�X�3B��U9����T��-b[���+i��3���eIq�ڊ�Q�Mc7���z��OrH4��nt�#���/\�h�u4�����^��9WJb���g��W�MK���mq.C��{�j<�X�8�/[��N|�*��hO�(G:5x=��}�t�-9@s~�R39�0l��L(�i��Rr\r�L���x�+|���l��Z�.IY@��W0\�"��0��kBmO_p�� 1��6�3�b�L�]����1�Y����tV���W/X�%	k�e;|O�@ގx�L�e��C"I��ɢX��	�� �����$���S��g��pY�#o�MJ73��"�Z��>�W��6F����Bh�mIOe\�w4j��'	�H�ܥI�hoia�D�ֈ��Y���.M�
O��x�䁞�["�W�?��sW_uY��K"H��C&-���n�����%=ǞMU�$�Iwm��3}]&#���.�A�U��4�;�����Dd��D\�C~��-��HffN!�s��URbk�w�����UzCW���d��a�LC"Է�?��S���k9g�W��n�$5�s��N�����!}�c�N���H+��ޗ`{+��R[���?�V�bg�J���H���V�ђA��m�Eu�G���(�Ĳ$�|����ّ#�X6�`�#�'g'!�C���8پ%��=v�a�g|��\ x<�~oMB�No�gQ�O��^�J���!#��Bn� 	0�_���<�ܵ"�߲����Í̐�t.#���Z��+����[I~,_����*���F�K�Jz��I�rAhm.�C%s�zm�'1�Z���g��K��z�C������]������>���BTtgʺ{�-L��0�%�ck��T%b�A�VOW�>�$��4I��5�Xp�{(��B��#I���n]�Pd�K<ޝ�C�+Ϝ	���� fV.+���'`�X�X$P)'u; 6;��R�6��@a>x��K�3)B�7S�F�[L�3K�jC��Uj<£�[8���p+�3b=b�xa#Dh�j'�5�o�ݿw>��PX���a<%���{�Pp;<��f9�0^"�}���Q	r��:����(��9���%�2��XmǝTrx1��\�Y��V.G�"@�G��&���&b�>���������O�ް&N��p"u�w���S0	�� K���>z�ў��&�	�N�c� ����SN@R�Ӳg�v{,.�͉�z%cvS5x;� ���;T0�Z!����Q��1,��gl��}=Q���i{|�~� G��9������ M���w�Z�#�j��M��8��8%Rژ���PkA��(��}�L;C�ܲq�K.�C�G�@s5bd�n����6���x�~��ٗ�f�uXlxV64EB    fa00    13c0��
Y
jF�~�G���i�ڟgPR緕�����g+��i"i��#���$�UA�ܰ��ɼ�U� �:�|`6�2�Fzv�QosIO��TݡQAI�W���Qq�oӡq��G3zb��%%,}]�)^��g<�4��fn��(�mA!������J�5-�?�x�̓*B�j�A��Cl��	D�U�2�4�F�i�C���Ֆ���(E��O�CX���&]��"��9�m[cN���K�Ş��EŦ�"�F���I��1�Q��j�Y�1jJn�t��/�:�J���U�-jG@k'��,�Q0���I��n��H#��mH�:�ݢY�?�]���W
aC�ڶ��>�%B�G�-���/t$��	2����B'��=���O��a��M ,K��O�������r<2�@;��<��ߎiz�
aGoD�Y�^ޘw�>�%R����G�X����]�n��%]�%T3����/�%" �����Y�<~ŭ�9���F}�, _����([��<9&�;�j�z�%��F�-������~i3���z(�ǽ����?����n�ެ���*�0�,����w`�g���Z���`v��Ξq��Z5�a�����B�����$^3"��o4]]��3*Ȓ��w��㞬f?la��l����el���WP����%�\ߣ�O�瓹�2�cc0��]Vg���&Z�vY\�����{Jt���.���:*>��=	Q��;B��q��?�L��c�7�lD�	:�+���lt�ݺ
�/٪'��̺�z�iK=t08S�Ǽ�PQ|�k'�'�eۈDvM�/�?�+o�~�#��n�?f��I /?7�bq�0��U(]��ǽ��>0�dg�Ԁ����ݝ�*(�q{L��EU���l��Ԟˊ�>���Jev�P��Q��E/��\j8�C�*�SL>/!�
=�������kcd6w�v����@���[9g�l�?`o��"՘�f[іE���}��������g��yg�e"��r)�te'�C&�g�*��2���c'���1�J�i�|I������<�D�Y�c�����9Y�n/G9-����y`�_��BZGY[�p�*��/����]h���Z�o	��B�%J�����
���G0 �b4�)s����X�Na5G�2q��V�����
�"u{د��OO��c��[�&�<�����x�~�F��]��Ng0؃D���gddW��@Q<�� 8�;�J稍�5�V|�����xr4;�v�D���O��! h|�O�C*2��
����_۬�(�'b~ �S֭l���j	�:�z�����B M%÷I�;�e����^��u����� ��VVT���]��J��3,���%�}�^�y?��>��~��َ�gL�]��m���ni�8�2� ���v;O���r�6$�� �z`|���l��wRC���G�Y0}��yٍr����|�'���z��
��]���v�5�NN��"����֛��`OP4��!��t�A�|s��R rn����GB��
8p߫.��9�m�e���qI	��s�LCj�c� ��=�s�G�p�>��EL~zNo;�:
8˙��U����K�R�ԭ-e>Z^!7=յ�"5��Jd:��P����(Hj�i�2�K��ò�c�O�숩��yؤ��=��hB�C�ޗ8Fh�5���'k���LB�^((�a:���?#��Kإ&�	{���&���S��g���9D��$ĩ/�Oj��#��ۭ�̘yl�1�����������H[��J����L.�Iξ�ȋ���n{΍7$o�#}���V�'�c�*Bμ)�1J�R�S��+��̎�oJ�,H��8����D�#���� �)C*�M��l�s��t�SU��@��K���6�.���Ϗ���dI��(P�u�u3V�<��jii�h�7}g7�{%��0����w��6�87<G5�����"�,��p���bOG�1��8�� Y����|LL���m�)�Y�u�9����v"���0�m�r�����x�A��h/��O�ю�,`<VzR�gҚ�
���5w&4el��	�:x��l��lto�p�"�o���K3�6����?���O.9J8[�!i�Kf�錊��44�:s�'%��~QJ�#����E*�	~F����F�Β>%XJC]���W^�Z
�M㙾-e���GLh!�5���h�� G{���~�O$c����t)��y{O�3���4jσ*m?�H�>a��H$B���M���!#5,�U�ߖ[j*	�dWu���p�D�T�G���o<�i�p��A��l�R��  e�ڮO��4�x�4���us���C�����RL���
�b�&���EN~���t&�;*0�	6x��l�nNa&���ΥE�s\�?�J��k�# on�㋵�}�C��d�?�P�(��^3���%� '�u(��V��%7��+�(,�J���w���H�$�H	�SX�vC/3"m�r�	�<�ۄ�j��#���"���ר�����nb!�laް8�E�^CB���<y�
?N����G7����i��+I�%���C(��_tg5�|���P�T�k��q	IG,���k�E��b.yޞR.��u�`S&&C`&����;BWW��Ҧz�^x��7��C�����Z�ن���r��rߞ���4�����zS��=o1�Fr� u W�G�J7{�BP"�wwҗv�rCT�Mȴ�tb�Iĵ?������/�њ���@b�#*�rw�&ʍH�R�;�M�Q�e�LZgo9	\"�[�)�1_F��tY�����(�xXM�z#�G��K��.�[�����?�� 4�؛P��Νr�#�!��`��s��dϐ9��0י�>��?�����T@�OZ����X^"D͙L��0����h�cz�W�$����8�_�Z��]��.�B��Ȩ*Љ�sQ���L�����I��.�Gb�I" �� �:���C�2q�����[�C�f/*B'���S�uW/��k)y�'�YM���7B*��K#�@;O�����0�b�����6�+�J��3��;%��3�ꙇ>Rkl���N���^PzxudsNnǙ�G<����-��༈�\&�����͖���	�m/�H�g��e�f�\��=w�4)Q`(4Z���wJ׼���w�e3��������e�~�v��WT՚+Y_�ɦ1?��U�B�he[qY��J-�����i�f_h�o�F�[��q�"������.�J�N{�<�5���ǈh�8�!�}G$�f���P�E�9C?F)��]ys�i���~�@��q���l�e�x��k�:���?�`ٚ_ "�C1vd�<9DS�fK��V�+ŗ�Ai�U��%�,˶�M�!�#<����x�ވAT��}�t��}O^�5�f&Eh�o>b���rX{�cն< �;���v�$U��͛R�>W/�l���d6�bs�"�
a�RJ0MJ�d>`5�8��4䲅h'e0��;�Y����z����k�b	'��%���%��Z�]�X�o�����Q�uC�G���� �g\�S�㰷��dL��	qnB�4�Pz��^�j-�6|gĂ媟g�,Fβ1�����ccmp�����O��n���#@��(y�+��>~��YRJ������y��Hf>�Gz�&�:��V���s�NLB����5z�kȤՒ	�	Q>�nG{w˪����������/�]���k�£2��&9�z����/*L�#?RB<0SX���n���w#bc��C��Wo�l�,|��&��+kݦs��I�
�(�� ֳD�N���j���u���G��yFi��4�)pL�8��}4ek���lY�`)ɬ$�A3
{t�r���fѳt��aQ%�`<���n��b�OU�[|&t�_j�e%�����#�/�@X�=�y1�.P6�A�
Id�,�݄r#p/������ى�`����ςs-�$6��b�Hw��� {�m�8��v���	�DY�ԝ��He��߭��VP��6�O���#(�@���S|X�,���S�X�ECX��ֿ�D^u81b�w�[M�#�"z�O2_��x�g�Vz��%��<�G��L!�:���â��y����*�إ��,�I���>��S���k��&����Tv��9:u�>s3F��Hl���A���)o$�_5����܃�y�/�O�ݳ�d;#(��7q�Vk4�EZ���6_ۉ�-CՓ���i9B��+y��OdM�_�Imh,���|B}����S������I�;cPJĚ�y@m�u�`J�5am�j�i�b{ܦ�Z骧���$=���A��.H�-��^^����2�����p"b���u(��3^�Rya�-�-�d_(�{ϽG)o>ܮ�N�`�"G���uYc��6�NzG�\�c�
D�"�̰�N����I]�W���9��N&M���s
���wB��:$��(��������i"zNt *����/	�"��^�T\��BW��?�B��X�]���Ӱ?(w�n��^4������t�4��S>��:�ړ�^zå��e�q��oH٣��7��Y��'�i�t���0�My���4���ю�-W��������]-�9	E]��e��.'��UYt-�'�ȪM�`�]�k<��&I|��wP��o�Mч"H�@��s��S����>���P=x�y�Q��hr�S<�Y3n1�]�mD�k��um1M[�z���a Q �q��}! �̌ʧ���6,���I����8C��(9�(��['~�V 떑`��7�V�3g�B��C�AwK���vc-�д���*8�侰))v.��ŒZ⢀��gv�d�7
�W�c����DCY�!BC�KI=���8�����Ί ف��y��ˏ�����g�XlxV64EB    fa00    1750��K�I[h)0�٩��|W���'c5pL���3g�8ϳ�3���˒�@�����;$�Ʒ���va�hw�O��E[�N3�5k�E�
y��0�"_^�g�<��
��Q[��x_�bˆ�t�	Bd��G��#}rS�����a��k��l �N�yA�$��݉/y��aw�fp��;ʣ�E1������g��K7�T�'Bյ�%�����P�L4��&��DT��w���4Xɹ�*�T�A"%�>��>� �
F�^���C �/� p����[������j�r��\��q�>7� ��8�:���16>	x��bA������r_"�1�לɸ���
8�����~u��m f�?���1��.�'�@�o�G�U�,
�2E02_� �)�?Z��7�3����a������ۧ�,v�mόJ�L�:�9��`� RV��8�X�sp��ӱ�6E�*���/���� AP�����)���k^o�V�6Agތ��S(��h�JKA�j�&"g&��h����/�����u���Օ���7�JHy��+|��`s:�MkVHK�zȍ5]�ǠXS6t�(�V�����#�utƑ(\�<�7��ʟ�`����v�?�m�H��X/Lk@��^/�[�	�T���D
�2���z��,�q�2���`$��Kar�hw��e�[�Y\A([�����E�� 6�8B��%�ece�#���I`2�v�*#�<6F&��$�,�A8��tP��ŷV�D�w揆���#>V��=�`��R�F�(7ȣÖ��~M$�oV���+��q�hnC|� �p.�D�JX8F�������F4H:�"��4� �x�Ěp��H֥|+zP�Ʌ��jk2$]��N*�Lmf.��B&���h�U��ԏ��OU@7{���}⎨aj~���?�
�����#NnZT:�ZCڹ�wC?��K0� tlן3g�R��iX^Ӱ��u�tS/bd)��磜��:�8���N5ˡ
��0*\o��4x�2h1x��;�ʏ�kXx���K�!��#z����w?�HW]�6w<yW�=�,(�3�P�SR=/ yT�2��q�$ER>�����!}]�OǊ�� ��q���L��i�,����eˑ���׎��w�{\��%9�m�o�ޒpH�(=��B@��hR �D�7d_�V�ʶ,S� e����T�"ߛ��&=�v�8!>g+��� ,�A����s^# ?�������<�β��_o�X�)���x��:�-�O�n%�E�g�-T�Qn�'�J
��s�S�����B����>xφR��4�2�v�K�XA�q�BY���n��: �+�������{ӵ��a��2��Y�7�X'Q�f<R��X��N�]��冸U��p�� v������eN��q�	t
�~��TA�i�_�S�� +�g��u��Ğ(��w�ϥ*���~J9�1��e�^)
�7Rģ.W�4�����/VZf@���\r�̼#ڍ�`��֟u�zd��@"&�M�/�{���Çyq��c�M����dbU��`�6�	/�y�6�6q����m��,(�%���4�Fg�!(�: �NO #�*�0��ÂHy��z�y��>a>���C��S��_��Ιs�A���n a;�o�}�SҘ�!�0Nx��(h��@��(�/��)%�Zo� �������n�'�˦&E��;���Z��4�3�BO�H���ShG��Ҭ�*c��w���E�M���G�C u�c(��<_%O9(�tOlƼ��<�ל�`��&������s�h9���'B	�t����v~�@��5�X�T*<W�%s̻U�N����Ch�����m��}�E�hrs�p����F��oP�'V�q�2�v�`��ڬG)�]͛���� ��(?b}�wn%ׄ�X�{��h"&�*;�1#�����=�<��/p��^{���t�F@�U��1A�%�k��Ol��ëDYUL!&	Z�+� ?��P�Re�]| �=\�ەl����I^97Z#���s�s��z�|pC�9�����)���IQWz:MR�V|v{��sG�� M{�F͇Ɔ�����vY��b�	e��s�@��):`D�;�
�M+���C'�)�1GU��8�x��9)!̔��҅�X�~ONI��dU��\����'y%�2�L龕�_�ä��j
��R����g6��^�a�~Wh����U�K��d"�<����1O��o���u}A����u�ų�9��q�[0�dKmT���y�F9��Fz�9�>qv�]p�>��3(^�z
%,!��?�+�S�G�}������� *�3��<3�;f-�
�8�u�yO����~���լ��"U��Bc]\��{�|Z۸�^́��PF���|��8Y�<����,��	���aaq�qC5��hS�+�9-jM��X^-����9%��<���b��^��g��gա]nΆ��2�B��[{P�V�A�*c�gaڊ�M�
MC�dg��ԢK��y���$#��K$��ë;��<�)ϻ�J����2'Z�^�BD���"|��c��k�\�a��%��<��hQ����F*ޑ�_����>%�Ϲ��#�����FJ6�S��D9�jm� /lV��E`E�#�����?t+�ęu�cp��L��=a�V�;����.�u�A���פL!��ٔ>9���5�
cW㙯�{�P�����#A�H7a�
��a�yYN��nW���&��uu"��@�]#I����g��Gv V��vQ7�}��԰O@���y�/.��q�y(L��ci����j��#g�ig�8FN_��AS���~���L���3uhip��E�0���!���_ϝ���s�M��{�!�B�) �ՠ���)R�Y5�~]>�@��a{UV�E��b
�JF�'hͩŢI�o�������[)\�)s0?U7/�'{7MsX( '��Fp���)�+�W�k�~2O(��`F�;��(���`���_�s�k�-����l�z�B#�|�駍��-�Q*�hM���^�o�Q$:�p\b X�Lo�m8������襯]��B9�0E��]���1������p�Z��.����q�/ͻi�#i.��i;��$s�S�7wB�!��H��{--;gŻ�k�r��}ҋP�&�E�5�{�1�f����� ���tt_�͆<�Ō]4 +�L�*&�\	^���^��O��M�;#���S��A",�#������*�<�n�a�W/�O��e�8�2�PhEp����6օ�ħ	q�D]��vv�USb��'����D��*���rV�17�x6���L�7�[�}{�B���߃�u�.Z���	D�)9�֟��CZx#f�G�1�PIO��9��TN��Y$.�c�ǉ$�zĀ�*@a����n�9�����j���=������1����BP���V2������UTC����gX��������)�Mc���3�����t` )��eϞ��j���:�AU-Y`r���Hc�XJ��7?N��;�"�˶M��f�Qw��P�E$QƈS�&Ke}���0H�;�@x����ۉ��j���ˉH���z���l���<o���֑,eN�Q3����VFz������8Ub���-�6���VX2 ��#��s�4����o����P�U��"��:[޳��>I��l�}=�	M�c�u�H�����Юp4��M��h����V~��(ڷR8���n�pL�{g~(�"�u��OHS���Z�ï��k�P4-bм�ypD[Gp�Z�87Tɴ�`{PĠ���5$���B�����kw���]Q[�/4q���p� 'W��Jǝv �;���8.y�
���h�V �-��K����jI�H�S.�|:��r�$˽k��M|�9�ى�b�{U��ͼ�E���`p�J���-tPz�ћd���@#Yc(-��<�y"B�Y�@��}/��K,�o����
�H*`�A�\�}�����F�`����s^|Kv�VJ"�q�W���Al�:�ķG��{�_Hɷ�q��n�1?WI��E��h!\� s�q `+g^�Qbdz̽����P\�2��%L
��q@�>�^�Xk�~�(F�p�����E���#�!e���9PMy�@*�~�/�$�	�l*���@�n<��|��#��ꣳ�o�vY����r�ȵZ��0"�^���-�փ�{n���n�otc�H���r}
�	!�����B��
L�D�i�乓1$����M�E���&�k�DSq�Zd;T ��![�.Uy:���y�"�L��_!����5�X<O�C���(��xp�J�FW�q�X�b"�גu@4�v�,v����t�(���\��@fD�'���}u)��K'�㯉�䌭|�
�q%˒p�f4�>Z���M@���ȧIH��Z�pm�J�Js��Bn�Q��q��ԁS�E���/�{sq-!��>	"b�KnX��k{���J���jͱ��1�_�}S3�L2��";���-�*�(�Z{�Pݷ}a� O���s#1t%n,�*��c6(G1�H�"�G��C�s�<Ҙ�d��t���/����A�S0�$rL�s���"7MMu5�6�MU���i�U��X���G	K��&PϜ��=
+�2���ƞZ0 <>�85�-���]�Z?��-`X�?���20�]��?�����brg�0+�7�?��Q�:S�.�)k�7;�s���{Np��x�i�l
ܐ�
��S(�Մ������wU%��@0힂"���UyP�݇�qL9?ͮ}�K�����!X?�=|���W��`DA����X��B���ŝ��HX}�	�����*b�>�����&^K����ؐWY��R��������[~��z;|`�/򹁕���-j��4�J�n�������+�Ĕ���Ɨ��e@�����_{O�D:�bXR0J�c�B-y�O!�%�V� -�<����f�(�i��c��������)��i�ԏ������O[��a���{�[L0Q��-�S#P�q\ /�1�D��&0�i��5��Y<���{�znAwg1𝗂����"p�Y6����νF���l�4�O�6j��$��9��ϛh�Rf�m�&n��$� ��j�Y] 3$+_Mͬ� ���)8Դ�Tå�,�K���~����T��B�����Q�I$��8�0&d.�?M�櫙"4C$�.a���XL�rW+�lM�ѡ�S(И%-�d���I�j�m�<X�Im�Z+a�б`b=�*_�7����N�N5n��
�I�oqch�{+j7	���ӽ��#'�=��g�ElR]�h����̤4���v��U>�4+���a�GO��C�%��ɪ��w�RJ~&�omxu�Q�瀕DKͧ�h&��M�=�������z�xwk6����ˑ�pj�/O/"�����J��8�`�=C	~y��L�%r�P5��`;Ӝ$t�m��GB����y=��PD.@ϝ���p�q6@|��`;15N��o�3`%r��d@!x��uu�H�Fǋx��i^�Deq�k[J5������ӄ�g��"�\,g�գ�Γ�t�]��ױ<��񛏛+�!M��{��§v�ٱ��FꗦR:�Z������E��V�����L;>%�������:Oh���!�Y��
t
�íEO���wAۓ�f^���I�>���%�3iVY�����	w���J�����L��N��p?��/�ܚ:A��T��#��HsJI0t�=���|����EK)���M�S�FE�o��)�d
T"H{������|����@:*@B�e�d$��򤰔�*I�;�����*��g/�4ϒ�`R��|1 ��l�Y�؆@�G���XlxV64EB    fa00    1840\�~G�
�y]��ZG1�9#�&��Vp~֗���}�GC��o�&����J4Nuu���I�=��>h�jS,��$+��Ǖ%x�ϭ�<��"g���!)ar��c)
K'E��� �U2�E��.��RP����h����ʹ��47���ߢ�wul�׳f���ZsJ��U1���ʇ%C���t��������Q7�W��:�w�s�7^Կ�s(<Ϳ�Y��g;:r:Ά	�B���䲲���wY�ù����������s�[�(ˏ�~[�e�-*��(�9�b�1y��]lŠ�s�(��Üv�n�UQq)3��X�����w
��x�j�Q�E����@W)�	��m��� �H^��n#���2LP�U��Yp�=�8�f%���>��W[�rB���i^/�yn��'����3�'�Ep�����8"D�]T#�b���vx���L���
{,����6ݪq+)��t, WW�ϫ�籽����c[��]�ȷH�+�|�^UL7�辽���9	#� 2����aM�P��LҢ�ֵ��oյv���c�oS�7KV}�~_�{]�ή=M:�gn3G�]��ll3��gdN8]�����\9C�B����D:8�{/��v�]�zSP���D��'/�c�KL��F?�h���Ƽ�&���(�,̣�����^)��A�=c�`�5�2�H0�ϖ{������F3���{�ڷ4���Ɵ�p��)�4o�_։C$�D���s�=e��j�t��P��N{�.k�&�mg�+�[��>��Q����媡�S���*	������,
|��A��ӳ;��+��-qE.]�yD��Ь?�}&vوa�/Տ�\��qC5ӵw2�bg��k����V4d�\x	��T~�� dw۠\1��2H����#�	S��}�KD��� q���"V��}=����%�5�(Ø��?��jn�Q�E�!��e���Ѱ�H�X��6:��O0^U�{eS� 9����)i���,�����۞�'�9#��Bd�P�	�#Up$�7"T�%��3�>�'�YsJ�KpZ�յ
Z�E�\;&�-i�|�\� ���	�� /H�o��^G"J����hutS�Zz?kP���9���9�-��3)��e�� ��#s���ɇl�?n�q�(qJċ�C���l�u�_�;w�Od�/������w&�\0?ڄ��R�Y�Y�`���J�rR}��E�9��.��n\�,rhr��0��\o!H5B�����m�$�n'����:�:��Cc�y���~��Q�F��[b����X?${���ڈza��4�	2���!���� ��C3���N���~�r���?���6�!�鐣�,'rt��H�����)4-��@A�H}C�H&ulQ�&��;�}�?�v�CC쬼��7�3�� p�m���~�"��V������P�7���s��ꑄ�Ú�I�
u9���52$1�� �����i�pY�^��I�tօi�ģqs&����s����;���*)ぶ>�`��X�#x�T�t���!���x�����V���!������,/{�X?R)ȏ��鱗5XiY�d�=�-Z��W|����0?�4��tt��3����K�o;BhG�'����,�K���{O�2 @�����5A��V(e4X�V*�+�֔�g*¢_{�=�����a:��UJ��]����	�H�r���O<k; �Д%�(^��c�H��_Q�7�績�_��{'6�`w���&�?�z�`�70�&��Ɲ,G�f����xB��&�`�>���XJ�O��,�,ʵͿ�p25�X��E��!�[�d���Z0��~��*��v7T�������;oyO���Fb�$������74�2=�� U#��^2��z>�Xq��G�zS��t$��F�FH�ܛ*P�O��
��64CLh�� !���,)��W�_
ud�-�%�����{v�7T�'6��a�	��`23x`�g��n���Us���-1������l�e��&]tu��C�^E������S��"�����Hrf���kJF�{�숤��mpK%Vp���� �Ծ�(>7�����/����}[80 �/ҕe[6W�$��� 3��%��*���j�䣄�T� Kۦv���Q݁ŒLuDU������Pْ�`���#ᰙ0:�S��2�"�j��r)�/�W�G�,��+K"$w1}(^`7��˸��M�0�@^kWB�߾��@�]��)�x`<J�s<�v�Ǿ�SsAyߝ�'�w����^�Wq�+�C�Ϸ�Ŗ��6Yy�&�U��;����ӷ+Q�-RC�yrK��k}�B. $�}DX��F������E+����dq��c��C"t���	7�wﶩ���;w�����lFZ��8�-.�E�R�۴[_�P� !��*&8��p�YI�R�r�<��>q��XS�vL����$(BK_,�!�'���l�$��2�8���r�Þ������S������pe�[3���8��7��	���|�X���V%�����_���*�rep(L.�~��M�*���qlB^�
�T���%���4@�cHf`<|��җC"Ͼ!�f�䨹2Ч�;NQtc�Bv�u\)g?I���x��p���G��a[��iTT�'l�oSn��������$Ɗ<��U�1rp�O�5d_�mH}���55E)$�^"�AzK��Q�`���z��u�Bޟw�9i������q�XP�~V:���+���)��v�����C��@�od�{^�mr۶z��h2�>(%D���9�Rݾfpmq~bV��������+���A���S���;&�@�p�rYj%m�ԩ��B����	J$ H币������(��5*�����t��N�8B�ä��)�@	�E��,�ڍȂN��E�q�Y��u�;���#��3��E|'���C\����$�vBF�;�a��/j��=��T!�������O5l��d�g}lW�%�s�m!�����q��(�]��Vlm���J�p��#V]���N�*m����p��olJ�3
���)�<��Zy��Uf�um�Y�e�3q�^���7�Ë�>C��3�R���4�yQ[�[���#v��w	�0)��.��^ȇ�+�l������ �C��}  ��|k�o�׿ē��TK�j��y��&����P���$O���G��X�E���	����̡�Nc@����=�3(�H�֓�^��<�!L7P$=�G��*����B4A��.�a���"��q1����J�T�#�3w�P�I��HmW��RQ�.x�_Ğ�h/�=�����c�����x���i ���=-)v��N�? x���M���?v�\�����o��p�Cŕ���m��>��s�;a��u}�=�A�N���.�� �a��\�%�X�j�i"�waӸk�AIDZHu�U1��Xe�d1�L�m�o��m:��� �� ���o	�wo���dWW�g�L�=���Ŧ]���Z�����zfq]�5n�v	�r�3گ�F��p�n��w7�8���qK�])�jtH*�3�)jV�%���o����5*|�#%���O�l����iz��y��R��aź��x>u��%^/�,G��8��ܪC �7�@�çL�ˎ}��ֆ�ͤ�m��j�	Z���!G6ee�G���}o�p<w҅�]	�	��Z�JO/��ë́�9}���9��K1_�@1#��&1��fJ�T��~s�ḗ6?"o�H��7��'>b��A��:�<;�+U�c(]�'��H�
"�I8H'6�ӿYeb-K��{�C�����@�h���a���kI�<,���vF�9��@��}`�����E���\�$��<�X:X���rAHG{	N#�-�8���Pcc6�,��8	.�v�D�W�S���,���X�C��}d8����^ȩ��rf�e��ғ���}:�B@�6!��\n����(�Dl��,wޕ�ܨ�1"���,�u�nm� &��:�ǈxk�]�-ZuK�~?��Ґ�ĥ��  �iK�W���Qz��n��{���ZI��P���v6+����7���̳&�8��a�t=�3>ŀ7�k�[<Y�Eǁ@Yx�8��@)c ����.�.�'��������,
[��$�
�k|X���^5��p�\�m�xgL91s�t�)O�쉖P\�P7�-w����y���8�)�x��Vtã�"�����.��<"��%>����Go����&m"�|�p��&���]A����e�br�R�k)�h"Q�UO`d4�A����L5���]jF_f�/{�Ǿ��4Ywc;)�5N(�Vb@rI�;"o�Q�d��D%&8�8��B'8-t�y�j�|�,'jI�ˈ5t{T�s{��L�{h�`�7^�`9�.�Kc�جFHx�z�L6>�
m�?�=��>�ϐ԰���`�DS�x�FY�B��pڐ4bXG+��c�9v�\�'�Ǻ~?�ާ��,�ɀbg�p����T82�|���3�0�Q�D| +\܏aW���}3�a*�̀d]?��f<t���l܆�?h�L����@Uq�����1�&������4���IU��N�r�V�D��%���>�8�$�Ća��^��iKi��h������%]k+����V�2�<D l�e���o&%Իp`܋x�IwnN��>�F;ס�^�����5�w��|�
&¾�� ��+ԅsϷ�3q� �s���%w��	xu����{�nwV'gM��/vl�>"ȏ��h�>���eP���Ȯ��4\Cy�V���=S�H2�j�>7=����v���}��F��"Y�����}��#�w e#�`h!���q$Wz�J@4�r�K�Y�[I���4������|����f]�$P� �U�A����~te+�3�m;z��H*'������7�6�Ж�<���(4��̂�u�������]_!w�F�q#�4t�Z�1���jA����:���#�A�vÔ�!x>��J�CU��X��0mo��*�� D+4�K�]�?{CҸ� 1�7��K,�qw�j�[�I 0g5"�q�Nq�oAR��Y8h᫡�hO��U�,�*�P���W�q��j�F�&i����j� ��F�E3̪��� ��U�r��%��};�����kتkk;~�����Ɣ� 2�W}���nv�l	ҕ$S�Yv�|shO,N��|gYA���qZɯVM,��a�c�R;u�^#���+��D0��G��MH&r�#��G<�wN�N����h��[�N�	;J�t��x�D�(R�~�@?u�/����&ƤxK�a�����|�i-]]�u��� a6���=�IG39��A� �ɋ�0��u/�T�*�w��PK�[�G�<��h�c��WB�ӇlS��}<|q�/�Ͱ0�������&���ޑ]�����.EsS��_݀*�a&䞭ҁ����O�Z��#ys�f*��v[?��'�;�z��=��$��(��S��p9���؍��Yf�v7�>��e�lc�����u;�<�.L4M���n�J�c��ו�����Y>��I[�y&���O/N25�a�k۱Q��4Wk���O|���/��Yx�NpΞ��lz&ёE�^�R_�i��r��pn7(>.
��Mj���F�	�+�لsz����N��B�}�%��i�h՚�U�X�X�'v���r�7x�l���*�v���Ѭ�eQu�� @ɤ�gF_S�n�ϞM�j��ިF���M����б���Me�g�ɻ�i��Ӹӂ�M��VG�)������t�׻y��kuN%�Ps`��R+�C�TN_�T:��a�8�{f�n��SfCo���-�h,�qǨ\{b&^����c�wj�:�<�x�'NۊԜ����3�K��"E��=�2��F����a�x�r�'D+�:�?�3�ʃ�c}F6���\P��h��e��h��^1��C,��ܽMF����S}3ɽG��P�@L��y{��p#�DU�4�`��cp�1����n���K�zGf{� 1E�D��[j0���F���1��V���w��hڦ�m��s+hK���^�mxK�9N��G6��=XlxV64EB    fa00    1210�CsA8�� ��u�F��M�|��$<2+���˵�O��F�/@���1�_����_��_kHK���!�K�ģG�י%�$>���*c��p7ك6~ۯ��7l�.��D��ٌ�+��QAD]��RN�4 x�샧��sp���l��#�1�g���d}(d4�L��j�^��k&&Y߁��%���c��U�P\�vj�ڕ-f�J��5�5�Z�v��'�<�Q,&�ƈp�8+��&��I�uě��)��U����3�[A}65�1��+�eq;NZb3|#].���1�IeV�aw��������Mo�e=叫��)�چB���6$��D��:rw2ԗ�oVB��7a���*ץ&��>���FNm�e�BH����MP��c���� ,\{4��MpL�������R��|�T��5���h�f<o��V�"�\&>��r����M�gZBb@�,��_q��n�0Wr�Ԡ`�[��rf�Lp]��&�[�w%(25�Lu4�Y*������3�
����.�(�7��98g�^N�G��D��H�����]��dVO��ѐ��^�EO���OͣS ���=$q��3���d�K�Ԥ5������["<0�{���}4X��s�~p�}�iQL��,UDQR�zo�����dF���2���f{���4�D���u�zХ�Z7,~K����
�GMX<��I�Nf���JV�u�������Йy+t�������%��Da#@���O*R��ޫ	���CV�Lf@C[t�I}�#M���R��ǮA 6r�!W�>��mE��̸����&�@�|5Ca"/��C켫)�<s5M�[I=ڀ�]���Z	/JD��w��kҋ:Q�¤'K��H4�S���MֶQ�ΜP�e?x�Y��S�rۘ~_c����ˢd# ԧ�e���
-��^�£ຒz���}jl�VP����9Xq���Vi�����d{�W^::�5Nʄ��0��E@B��ƚ����6�� �p��`I���>rW�u�?v~%�4Wq�=
� �%x�guz��e��c������������5B+��z���@��sd*�0r���?N��_��.h��A��w�ȵ����c@y�{�	ƺeФF��º��Lw?:� H��3W��=q¶�Q�$�mp��%X���)G�|���P���D��7�ل��"���9l�SL�c��4�r}�sݖEO�F?�Pb����ҽHs�~k�L�g�dҋ�o�����SZ�����EC�qM�teC��14#�x���e}����X���dC� wC�v����90�8E��^ �Pq��]�qf|�4�����7#-�7����o��Ɓ""*َ�&�Ǽ�f\Ƚ/xF���d0W!��U�>�jh�����d���ϭu�`��\.��ZLb
,P4dAGj$�[�,7�Y+�O�F�ta7 ����r��Ճ]4��<�UΫY^�*Mۑ\�u5y��z �6-'�uC8�U�j���#�p�Z��T����Ŵ�n�k�r\�(΋oY��Ů�<�F��W]Ц����w�Kz�A	,<Z��f��hR~�-+G0T�8��؁d�e�ԐL7k����5^��O?���,���JNe1߼��$�32�D5Vz���`���t��grˣ����<;����ٔ����l����E���*���§��?�/�T,� ��v\�v�ăh#>˾��@�5�N�&b�2(-��}�8�:��7��O35R�7�7Tr�`�^��!�/��Jtm�s��}�����C���1�"l�u�<�_�^���W4�sq��5z{$GQ8dM�];�� �ه(��R4��x�>j��\���E��^�����fy�%�����@�J�"N2��%az��J)���Q�O;��Ԗ��,��ryp��?hَ���bZW�4ڀ���RHgCP�l��i*����"�e��W�,;b�-�t��`DlƕZ0kZ�׌g`4�[&�ȵ/2o�d�G�b�9�J!�c?�\�Em6sOT���T���� �I-ۻ���Z�'��1/tP��P`�~��9�b�o��p_E�
g��M�Z'�-�!��*��,{��e)���ѿ͈�����(�����36�X/�
Y�M5�����؏~���)��U	� ���Ǧ.J���>��n��Ë��4�B,��c}�� w��,A\K�F8��ؚ�c�ͷܥ'�����[Hj#�o�w_'��+�I�o�H�-�.k� ��լ� 7T_�L��4�w���WHg�����CB��M�������Ŀ]�����G�P��*����]7�X�ChZ���2nIO'-���}��5��&Ā{I놕�4t�V�����Q~� /ep��N�|�=����C�W���$�a��BUFFK5LLo{ԺHm���A��C՞�DPHܮ_Arw��-o�ߺ|8u�`���ƝM��8𫣋\�mư���ۛ�bǉs@�M���L�,�B|����x�[u���u���D!�aA�0 u;��A�q���� Jh�׷�,/I
.������Z�>�﯁AS_��E;H)oG��	��'�Xy�֔ANx�C����I���5�ׅs���������*�C���|v�����bYj�pVI�Ro����¬P a�@������5+8�C� �2��u���@�&�8��%���f�R5(N5@ 5�omBl�=4`�T�[���;	����&��M�w��HD�0V�����0٠=T$���2l���R�v<�ȧ.�wg�h�Mޝ�Ԣ����M���7���-h�!����BV��AY�M����0�V��g2�X�./w�!*�R[���,�&\���3`�@6�8>?.��/�(B\!¹���O�j��yq`.פR�(�+uOLC{@oc���D�BZH4�^�����פu��b�=˦Ij�g�+֫i��@�G�`��a&� 4�<b_�xԱP+>؉�?=`�0�J;;rH <�(������`a��͓�����t�Y����%gڂ/Q�;�Q��J���]�o �Q3��B5O<є
[����rHg��^�1 ��r=Η�m���t�k��Z���VG[�{,�X����M�L/�/�ڞp�u�.�s��ҝ������<ldNQ)��g�2�7��q5ɳ�,E��I���D�2���t!���j؞�����ҷ����ADe���^�����J�ˀ�{��=�B��ϡP�Y#^�Po�Vt��x�̩h��y���ɷoɗl��U�ޮ��|w 5��U};~�^���jG��)Uv�[4���R��1o�c���ܟS�I�_Q�����cp��w�ǒ�t��=�&*XX� ������Ψzj�V<`w�[�;����_HXp�Ĵ�k?��I@�e�V�U�~?.���m���V�pP��ʆ��,	�-�_p;�O��%�)�
L�irľ>E��db�$�0�"���*s�Ü��I1���\���姦��%���)^3�wO�@a�@*r�qX�ļ���"���'z��^?ԖfH���bam��;�����x'PB�(B�A!;�.=��)�{�4�8�Ã<=o���F��+3�_q������:���sW��_�q�c�êKw86�׺F�5��i�,kAd�T�un�r�3�R��"���7%�;�X;��{]QS���c��U�t���� ��7������T��-��.�=��+i���t@,p�/p��Ep��{��/�2�ߜ���K\�ٯ�oW����~8yz�pT��*1S�"(��:=��X���c; q��8yܨ�i{�/Ǒ����ZkT��q�ژ��[�D�IU����.$߱�`.�m����<��Bj���A>FD?���"�o�y��V<0�>�	� &+v���y	G�6�{S��p[3#@X�Qx�|��_�<�}|�i�e��e�G���~�!`�+J�Ӂ��h���U�p������G�H���^WYO`����V,��۰�@e����0�ۈ�J�.q���������i��e��ܠ���v������s��q���>E6��ֲ�DH'����M���L���3�`:�*�`�xI�� 9݅�@ �Zw�kzpk�ґ�X��x�8k�_y� ���1+���$��+|��Q=v�dy�N߬�`��@��W�T�$<���F��*�.�=_�><� ����]�Ԃn��*L9��̩��ctqPe�4�V�c�Jq&�oW/���H�fLƔ�����/SG������6�O�$Z^ab���I/��u\��9`J���ݐ�ʕ������U�e�r�"��)K���q�75��̰��bQuxr�%T���������R�߇syR��V^%]J^�w���K/&X��hac�Mڶ�~�脼Hj��QS�(�ֵ������[�wx��h2�7YQ{ ��ۨ��x�0v'�ҸL"����^+��� -c~k8�#q����m�Ρ���:a?���`6��fْ8L����i	��-��5�/���N3Z���nI�{\�֞y�L�3]�iXlxV64EB    942a     af0�j䐕��_�����r��Gb�[9�r�&���h��S�>8V��7��v�%ٿ� ���?� c	89��5�87>�r��/v>M�#����gX��l$~�61�A>����!s�-A�+o����I��>��V]h�xK~P���x�T�ܐ�+3��e���ܐ��OH��+;��͍����!��0����sn��B
�^<~�I0�5� �zg�J��d���v�yO4ʔZ�*�s,Zh�zN��oL�+�*������{ z]h�bV@��n��K(,�F0�j�%�Ũ���>)����k�[%�ڥf�oӡ��#�`_�~���{�Qؿԕ�W� ጚx�Y�`xL��{6!?����~����yyj��c�ڗsOq�6y�j�n���Js��8<���Y�s\<�k˒��µ,�k-��|�YH�A��K���O����&����z����b6.Ғ>�ʴnGɣvi�0eG���?[ëtZ��i�т�C�x�/��{��v	�ҟ�[�:h��ʨ�ʖ��~Q}3������{E��������p��R�/^�K�OA:�犏Jۢ~�紎-ZV6T8c*�08���K�w�u�&�7��N�@}��3�[��^|�����p�^��ba?:/�0��t��>+�"
Lկ9Z��g�.�V�Bt��qU���E�]�m�~��B�A�7�Ok!ķkP@
�z���_�l��{�
װ�y��/"t���PJ��Y{��3M�w�3UUTXˤ/��`Er-��A�<������G>0����7i&'�23X-��S't����z����5���lr������ll8o��i�51�ɲ��S����{�A`G���9\�k�#Y����~��i�D��8K°w>��n���.�Cs�/��R��Ѐ�S�ɻE%A��I
�����˪���qO�qm��ya�9�w]�s �Q|`kU2kzG��,�?�m�V<FR[�S�	�ď!8�xn�1��ح��$sCO;�]L�
Me�X�[�y%d}k�����PE�K@5��iz�B��ΆT�&��m�'�&2�����Z[�LȭK\H�touZf�־!�6ݵ�ߵPc҄�0�y�R�ѿ�b���|��Cx�ջ�FjC�LJ{m���5�G\E��"�r�b~c%d�}S�<�����O�%�'n��f��T�A�N.���m�:1 _ �
�hHl�ʻ�Ἦ3���e�M����M�c&��P���#��b��E�r�曱eLH�+��e���=�17��L��G��Q��� 	|�[M(o;
��r��f:�����w��k�`���W'��jڈbl���B�Q�����)H�K���~�D��s���Bћ��Z��]z�|8�3�!�F{�����i'�0��Sa�i��f,�>�ޜ�CkTs��Z�?z�4�V5Z7ڡ�E��xwuZ{��]�6�o��M��||�߹�3$���
A]���߇�sL�� ��[��4��Ґ;ڡ!E��bAg���xt	��P�דC�I�ȶ3"�k��t�gRA��/�d�L�e�M/�9�)B˔������]b���ذ;��V�N�z�#Hd9"��x���H��%1n��ܔ��F��z�ܓ���O�Yá0�͛�$Z�9��7����5��H��d�=��Y�;�)�P�L�E�ā���:�����u��0,����M���W�ޣ���-�~&n�lK9���Ӭr	����2L�c��s-���s�):���r�{O~ǯM��-p�7XQc��$F�c�ˢZ]��/��i��a�%bv%F�Dq�5�`R��[V���V�T���`�9����LG�TM����������*�R)�8��P�� ����l#��D�@ �o�o↚�#�u�ߒ�Yy2@rt��^�ЇmT���Cgl$Z�-y�δ��/�GKg���qi�؇b�i��-�3+�aUJ��/�.5���^�Ϥ�K�B�f��qL����3�� R!�2w�W�yfEi/��
}�#�R����E�8�
��5���h?�����:�����}��k#B���/�!�N&NǱ<�@�9�6���9�"��;���Wަ�'L��A��L5�~�s���i<7�B�G,���Չ�$(\�@lG�,1�b�Dj �pRՓ?��C�F�<ˏd�)��b�(ê
�1���܉b�%�f 3����+y{z\���-��y��S��dN����I-�RQ�^�m baq��O�ޕ'��P�%�~̔���7�:���#ay�ݦ�`���B$I%�ѧ{��X�4킟�~���|V��6H�a���G�j����?�Á��o��я�Zh�y�@� mQn��ԄP1+o���U����j��@],h���NL�LĂ.� ��B�Y����
Ụ̋���0�>i�ԯ0m",��VE�Ý�M`���E��%���e�VQz̾�"P1�e���B�����ӢAG��Ҥ��A�����P��q�4�{�^F�� ������t\zf��1��FFo�{M�q<dls>e�S-�.��s�+qAu��#����M����V��⁃x�3�Z8�c����9r��<Ϯ��?�q9_�N,�K���yo�Du�Zeɔc����+9)$�O�&>�8�W���)�ʯ���
�?��罋۵#�΀R�����^�+M*3;�ć8�DIlЋC�&�些�j+7ǯ::���,;���z�"�}8��_Sr�c�D�"�T�uR��`�&�*19���)��l�?8G$�������g� ���{أ	