XlxV64EB    1cb5     940�m#T Q=_�u
�EV��C�D��;ף_{_�^��ʁ�Y�:U0��UZ�v�㶈I��6-��J]ʩ+�G���áx2��>��ƴ��8�w�,�5�[g~��N���d��R|eT�R�.�(�O�f�~C��㫖oC�^�쇿aE��-\~C�y�6]̶��n!���,A3a�(�e���MZs���c�R��/,\��7�e��ͷZQOV�ȏ.<*XA��G�UZ�Vh�@�=kx���tUZ$��G�Y��Qpj�'zHп(�� T�"� ���@	yD�84��>�֢@���P"-j� �3�{��Lׁ!�o���[EJd�z�c+S�}��FO-���f�fEl��^���҆$o��'H���%p ?��L��UƎ\.��6����k�UՇi���oIzMo׈�؎�a������.c�_�o�CݖH��8��ra��&���m�Xh&���5�I۟�p�7tag�`z��s濰�bY�������׼��X��A���Kg�'���U_���N�6�͗G
0�����<[�G�D�L��M��֖M��m{kgp�/K������k�����T���>�sJ���0{U��~��c��T<@�-C�H3�9��F��I\�b��((s�<P�̊���:	�7F��-B�s]k�>�`�oLʔ#�P����J���I�kiz1g],b��ڃ2�;?&���p����ЁN*�����y�sPY��?,P��٤�4؃^(}�Xk��P��/  ��}���#�U�l���4ɔ����6`�q��R�2������=�?tŹ��Ja��^詀��̿탞ؐd�-�p5.�,�5"�K�D=N¼�=����-�E�ܑbL8��V|Xg,:EH�<Rhɥ�*lM��C�]$Bw���-��cʺn�I��0��W)��`�~���-V[�P6e:7���E�ǫ�����@���t���T<�)���.��=ޟ"y?�E����������N2��VP�`o������ ��mzy��C�^�.F���]Ż`?�]�ePE���;*�Ɖ�����g1����wv���Z�?Ң�hW�����UM�$~(�J�]��e����$�ٶC�x�< ��])���4�¼�x{Q+iNWт_f��g���>�9D�y����,��+Ƃ�4j�sץ ����%���3v���i�6���h`�5���o~w�MR�܀�@/�7�%&w��>,_1n�hO|��,3z�*LZ��ဘ����J����%GDsS�K������|i���+l�~�-�PÛ2�ֽ��\�m��Q�-���������y����h�1V�1ZD:��l�8�98�O�Y/L+#���~3��g��J=�zrH�Π���,��|�~mV����th��3MXU+qî������"B��}t���!��Y.�x�#U_"�.�F��l���GC5s�\��"N4z>�fY��]<�֡�܎c������}�3�;��[�K6�q����)�t��D���a�R�v��_l(�F��Q��@=��'tK�V��P�=bs>:��������_�{םm��=s%C!h�5�L�����G�n
7=u���t��q�s�Ƌ���`옺7�)v#X-<�I�q?[��J�-�4y��X��ǾF-���ج�J�yp����d38�e����-x��3|\Ri��1غP��u���Q���g�`�.���i��O3,��Jh@�;��Q�h�����������\�]�q'���J,���h�5!$g���Sp�%{��~f�X,���?9$g�pC�S)IF:.T��N�O�4e�h��|=�9�3�E˕�l�ɜBI-�R�g�Y�"%�n떜�'.�儽 �6H��_��4Ot�l|f>�̓��b*���u^��~�����������B�"OИ�]�A����A	��kD���	����u0��Ӷa8 ��*t������QE�����P�l�=��v8�7�ƃ���M�1^��A�O(����[X��g�6��>:���_1���Gy�!b��Z"�����¨����\�Rʲ%O<�6r���ޖDgIY��]T������
��8r�7I�����$�,D+y�ok$D�ik E.���Gsd�T��P'�Y��*UKf*��!S�̂�[�\���)z�0U��׎d,�>�y=9���G�Z��9I�2��?# ��# �}"q>��g��*�)���j3�_�f#�:�>۫�2˺^�R�[R�r�����c��<}'p�׷�M�vB�������BѮ��E#G<,��Z�