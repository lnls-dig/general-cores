XlxV64EB    182f     8e0s�#�rϨ�`P�bwKv��?����Ӝ���Ge\9��M`���s�}��C������o>�e�}}2�}���R�c4J'�g��䱴�������ؤw"�H7������Һ�K�����w�w���i�^C���{�,������Iu! 6�>HA��Z�q�:5+���{���	����*\��V���t5���oG�FF� �W�'��}���?f!+�'�ʙ�yd��I�JyF�Cv2�>���'ϑ��=��d�	:���ʕ�l�E<Ӝ:�.��s�F%9PQ�m���Q��D���kO����>q�F3(�zy� ���ڽ�;%9$Y���6�����ze�ܩoZT�g�`�D�����vI���0c:���,�h`�^��ur�1 sͳ����R��Øi K>{����2)�5!��׋H�`�gN6r�����ر�1c�F�b����[�Vr�OX���m'b�nx�P�/�]����`�@�ꆌk�`�9�<�؍�XzL���oz�7J:�ح�@������^�ڴa�Y��؈8+mB����1�❜�t�Tb�d5�Ft`*�Ng�sڥ��7��#��a�c,%��ɚM�G�����D�$�""��R� F�];ήxb�$^����u�����~>`m��/7ҍ��:`\��ΤD<�����>��':��ע�5��C�>��_gM��Ixۃ���j�E�x)?�ޯ��0��|	������}�V�	`��gl6c�4�N�B�/�|<��#�J��g��b�����Z���^I�'�g�g܏�NI��8�*��E�U��ן<ʃ�O�CX������R��W)y��D��(��x� `h�p���sp,մ�(<s�]�������O="-�!*�IG��)T'��wh��4%a�'N �,a�P9�^�OQE��|�s},�I��O#HP�Id~�k��lY�,��]������4*��M����p�b_9Y�fo�̊��a"e�~����Wn�w��^*1|CxU��b�6a#��e]<��4�ƃ�:�Y�"�S�T�_����S'���ȗ�c�{��
�L�;e�Ǹ#��bp�n���~�}�D�N���R;	��Y�GI�
�?!�w#pJ=�\����<pu\TL4T�b+Z���Q���,Ǒ�GJ�$�zk~��镟�b��pvy@���I-�sr��s��_��s��u����$9+>����-�6
����aA�dV�l,����M�f1Gj@�x��W�]��*A|� 铡\������}x�A�B�pp;����+1Ԇ�ʋvښ�V�[��;V�
�M8rf�:Z�5��]���V���l��TY�jlص��C��#�����r�ݧC-ˤ�n&��W	,��W��`,l�Q��F]����N+���3m�V����TuH��� ���?�n.%>� �5�5u�~���w�V�o�s��,Zᇱԡ#-ɀ"p��_���m��˕�t��8���׹��:@ey��y��-��/fB��2�B�D6��3�_�-;Я��_ ��PcF�F�:���]+N�Ob#i3SJ׌-�3�8d�ZB��Sl�����4�z����OB�x��u�wJH�oC�W�}h@�"��B���E�+=�=�ٿ��t-w��=�e�K�Z�<|�PD�M�g��lj��|�cs&��(��d��1����޻&_QVրk
!��e������P#��a�,�g��x(e�)��O^��)SB���e2��P4���m�t��U��WV��h��:����j�;Zv+j҂�&v���b�#�z��o& z\��������G����N��z�:�s���t�s
$/���P~yHZ^�ڢ;k��&A���L	�}_��s)�uBO)�]@ Z�ter��t/�
�]ȭ[��KG��Ϝ��&p������*�`3�����"���<6],@r���ހt��IQ�m�Y�طy�8�PX^��!�A�����x�4��X�\ˁ����zl���]��{�v(�	��vpe�>y��rY���>�6|`S��U��$�z	�۰�QB=a�r���q��(f81!t �?���"��R��|�r��w���zb;	�C� �Z�<{#�WRĵ�	���U�C��D��HZ��w�d��ߡ0/��V�h\Pb���`6�{�"8�����F��1F�<�h��0n0��f�"�z�dz��e���}�]�j�