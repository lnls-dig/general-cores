XlxV64EB    6378    13009jb�����yy��ncG�R�h���y�z�L�:>��������K�bLU���E��7Ģ�@kϿ(y��Gb	�lz_ �Uee/��޽�%�$M��Y����(}B��^x����$��-*X�[ l	����8Ǌl���A	��kz�o-��j#*�z���zL_Qn5|dj����7�������`���lh~�zډ9i0_>�x��C��5��WP4L��/��u�K-�=	��1N�YP���u�V:�~V��}�c?
���rv�ECĚJ�~fuV�Pr�{s�Ӱ�i���(�S�1%Dи֓*��3/��f���w(�wۯ<�mw��QQ�9�Uz�q��:�߾i��DO =�=қ�I���p�,����$�P��?��蘨0!x{���\8���(&��fs���۰l��Vfc�A;s$�wc�(M{/P���h�hR6\� ��\�A��KJ>�Ǐ�ґJ�*����霤@x���d�E7����;�E�xF�T�p!���㦺�� BgC���/������ z�U`۞��X��i�5N�1Ō�R���.�B��k����� �c�eu[K�5��F���J�o��Q�?�|=�ݐ�;�xc���SՀ���,wxvd
kƨi���m��u;p?��h��Uo��/���C����A�Ǭ��7��[A\�m�k)D�xo��KX�Ǆy:����J6
��U�i�ث"�$;��~/���w�8���0c��19v�WZxI
��♱iR���T�t:�����!�A0{��f���xH�er�A����LoSC{uE��h��c�������J[~�2v��[tERc}�ȪҘ�'U'M�f�q��~ѷ�&Zc"9�;�[yXػgY�d(�nB��W�0P/��8k.�7Ԟ�aO|���@,�<�����^��ED��{��7���6\x�@�\AB�T�̢?���ٙ�ۍ��A)�g}��=ul/�ͺ$ژ�\ӊ�t:8�[L��	~ԺkK�T�0�7.}�b�C��7D4�8v_�X�
A�If�D�>�U�F��Z�-���z�]V��s�˾��2���Aa�_O��I�k��H-�34�q˰H'�]������?��h��!_��?�n�t��%G��k���b�2I�E^`�Q��oi��)��� D��Ґo�� ���g��x�(9~���cȻG�iKa����{gl7�Ƌ� _I��u���k,�q)���"]���?'̓0�@�����	�3)�w[Σ2k�jP8�-'�)��AN�%ke47$�<Q�Dpf���g��o�FC�b����6����$���-k�Ke�1k���I��W���j�E��C�>�j6<r:��ۭ��V��;�D�������WY���D���'�S�����ĉ�M����z�d턨Ad��ƪ�� �s���N������ђ��T�F]���ы�[`����N��zſ�1��E�o�^�w��Q��|�ȕjS8�0�:����P��=s����F���Q��w	7�䤽L�� �O%v)v��	��H +;(�"�r�915*��Ͳ�;�b��������jءԐލ��!���TH�/TB;v�R��K�x��:���Lo $���+k��9����$�G�x ��l%+� oR��8���%S��eG��8[?��e�S�S�� ��d�?(�lq�Q%�4ͭ�J1)������/�'�͓0��p�h�M-k�!��I�s64m�W�/�4u;PGv��I�AȌ5�SQ���7�0���fD�o�-(�c�{ఌ�u��?����(�反�e���ɫ?;(��<XY8W0b����/�X��Ȝ
D����M�c\�zo1�CA�� �����L6��y֬�+� � m�)n�J{��I�A��X�������b&׽�Bg���	�����+p|�/�g`CgQhH�C8D6�{b�iG�"HY�GKu}4�A�/\PD�@����f��D�6�4��Π��s��;-�_�Lsj�uY�.��j.�M��v�Y
��2�w�m�č�DSQ���uW�~�Y�,�+�`t�D��=��Oq�PkiX�6����~�]/G��V���e��3"���-v�6�E�"�o�� ��Y�w��f��E�:����������`���V���m�?�sBm���Q���-�S��Vcl�Pl\�`�u%z���o���'�r_ʄ�Z�[Q���7g:7G�mx������V�����"���E{�-3�G���O�_�!+���q�gMF4�
L@�tf�:���Lε��*�v��>s�ݽ�x�H����샋j�B�*�����nۭ�yFؤݨ:A�{��
k���}K/��_'1&�_P�c�ȸt��c�j3r8y"�w��E󻃍�����U�Q��c�&�U�ۘO�{�d�!��/�d�E�bZ?S��c�٦
:�9�ݢ�f���Q��r��T�`'���M,1�;�3^\V���J���3���邎}T91���V56�������4u�=�&t�h�u�.T�OP��U�>1�on�͙�CNJ�`��1`'�=�.P�Ks��>$k�2�vbTp�CL ��A)�eĎ�9\
/���g�frf9@�w�_���@Qf~�raG%��I��#P����������W�X<�I�.��p~?���/,;nL�
C�Mtf�1�4�)m{�Y�Z���cf����[Z,J9iA�l�9^�#^���NY�� �2����+����0$&���z���N����T���&I8i��ZÞ��>p@U����i٩�3��A@yZ�����`F<��8��# Z�y�3�����h.�4���z�=�Oȶ��L����ޅ�H���D��x5!��y���}����f.�P���7���[vt�X*3�x�	�,��(��3�T���Sl3A&��I��R����3���1�ޑ��ڞ���#F����K�=*8���7���\���C��l�w3�C�{� ٟf�F�/�ˡU�$�Ty�瞄�Rt��>�P(�������F�_�!z�!����eɻ��ô%�D�[dՄ/���2Ὸ_̣�qm�8*X;�X�zC�{��{e��Nom�Kl\�8�ыD����{P���3J�侶��~��\���n�K}��L�o�C_�װ��;�]7*e���E�dT<���G�����8:%���&-`}��E���''5�������F��h6J�FY�����/]�{�����"����/�~�ۣ]�hcYwڗ�vR��ˣ[�����gm��*��7mr�Y��+���d�A��/ �0^��#��1B�k¹����ī�/z㶛��_�>]��xE�@i��P���iڧ���v�`e.i��	��Gy��h�s��H1�7������J�"���/���_�Ǿf�{s6���Q�d7�uF5�9�o����K��V����j$��!�^6�'.�'FD%g���ηғ�E��l�H)�Gau<�����ˎ\O�Ҁ�	A,�t��%vt�#��r�H��W%���cVVF�,���lm���P��/���#(Vf̠��/pj��$���I���Z)&��{D�e�(G�j�����R\ܽ��՟��F	��?�t�����Ə�,���e�)thj>Lm`������u,j��FgE�$��jAVV�#	��I '���+�K��Js�!�Sֹ��l�jCP�i̲�G��X���1���g��S�F&�3��v�Cf�qnY{����~=`�H�!-e��CPX�r�/�4Y����Q�:e������	лQ���Ë�o�i�m��x8���f�t�g-�ͩ��Jȝ���^d��O�K�b&���O-������0��nֲȲ�j�5�@<)(1:b��y-��o�M�e\T���1������o�;�p�D2�rc�D���E����V&żi�Na��Yt��Dap���x6������A�~�ޅH.¬�-��/7hv.�Y ~���h��x�엡��뽟���Cd��8L f�j 	 2{���&L�Lo�k5T6�W�'�D��5�N���_�>Fa��Q&&2���6��4g�I�,e�{4�?r��7*=i�\�A��_�n����tw�nt�Uï|�Ș��#�k}=�����oE���}77�f5�WM�&uS�Vh[��͍�3��DO�G`ȻB��������;�sC'�m|W��i���B�	�wG��
���BJ���s�V�Pצ�e9��{�n���C��6����[�<����v��'��	�Y���%#:}�Tn<�"�R��RRZ��Y��cd�^c��?I4K={7�Oz� �mNe�l�-��$�I܅���{�-s_ ����2��)�j�1�^��"����� ���E����)�o�>� #}�,q�j�9ށ�D�sP���5p��t9���n��ck�7�͓�V�8�d
�<�qѼ�ƹ$j���G����Ǎ����� �YR�XM���b��2�Q�Ǳ��Htv�5�a�Xz����5㲜c���k\��B�[�R�⹕���8��q��������9f����lBrI� 4LkE9 ίA�G�+8�9w3�JF����G��ru�5���]iŸ]ܾX��எPե��ψ�]�b�tM��ϱ�q[̶G�6���lx�E�0Ȩ��KeY���W�g&���z��״%����e�n���z;Էkc��r�3h8j��P�H��REq���]�