entity xilinx_dummy_sim is

end xilinx_dummy_sim;