XlxV64EB    13e3     790A�Z��^�Ə��М4Z�a�V}ɖt'$�.�_�]f���~!5@gu%�䔪 1#r ��A�4�,6�#d�e[� ��k���^�U������b��ٱ��!��@L���q�Dj��4��
��
�R�	ȱ>�O�J�b�*k��p��<�Q�1�C�v̖�x`Ԝ�9�(�����~J�/aP�hN%r-��ӋL��r����C�_Wt|�ܫ�B���9�&J�x`��+}T�̾��ɨ
4�e�S��_:�
�`Ҏ��F�j�
N�����j�j��u�do1�((&Kq6w��ߗ��0l��ö�w�h����%���M�k�1�-��k�aUs����J��g(��ѹ'0�kL1S�w����X�B��
�x�4���*���K�<x�ipm�>QI�����Í��{�.!�-�s���/7�|4���
� |��_���/BT"@Gx�L�]��e�\V�Yd��=��O�/C�p�J������ϡd�v���+Xxk�|��3z&&����=���/Q���pwFD�{<K�л%�o��k"#31�s���l9�<����{�����e�q͒lFv��1BR��D���ǂ�@���r%��z|��ģ��a�M�F|p۰�'��R��T��cnz)�+�d<è���ф�eM�FTJ�1�[Yqg!XR��%S޴;|SK���*���׸��N";X荭�߻D��_���(l[�k�!
�akh>AK�8�l��L�Vy81�§>."~�y��*��J��%��E�#�7�d��P�@��3�y�M>A��E�i�:�~�>G���S�ګx�ԓN�ji�I4�7Ɏ���j"*^3S��Ԕr&��3���@����|N���ӌGR���<U\䘕���bU|ыof]�� �onO�>��d� �ٗ��,����-l?"�ۮ�n�h���p�Jk�95:�����͏�ӆG�]U��1�F}�ok{kj�*�h0v�\^����)���=�3���oP!�О��<ʈt�Ӊ*����-U$���J�Sr'��	�"�Ԥ_n+߅,F����r:��}B�-��7��%�2���v[��*G��dnU��
�Q�@̗Ȅށ�!����}kN��{���Q��_O������V2	�!5ꇰ�,,�I`��ܗՊ"lK�L�O� �:� '�Z���X�w��_��}� p�H��ݐ���㏄����,�i-tM��i6�SbP�ںTct�_��I(�ȆI�`����/�[\�w�
���ϣ2���Bӯ5��6�Cdfv�l	�-+<B�n��n�KY���RuD�eL�C��{+S�I,ƾ�5�g�a|�ə$IMih+%�ُB�j�$��M�uk�wB]ۥu�"��;�	�J�~)�s����S�ʿ��r�qM��Fն���T�,&NeR���$�W=�?'#l�Dj��%c�G1�j������@M��M�]&F�U-H����3ԇ�
̝ V��Aq�!�Ty;H�?��yGE�I��Y[���'c�S�,�������Ë�b;���Gh �I����WF��/M\���������1����X��.Ii���/���\�9��O���y��3�&'k��Ū���?��v����+�==:I?]2
+�d���>�KFf��~8X����:H��z��Rmsѕ�oTx;����b�.��H���F�v=�����o�,��ͦ��dL�%p�1�pi1B�j�h���Bb�&I���9u��p��p9vh�+TM#&U/T�	n�b�R���6I����M��~� tq�l�y��=��XR��PC��HuEt�{����/��X�]_����|xu6|v��N�tS��_C(gQ�J.��'��(q�Q��������i�C�'9ѭ��FUA7TZ5Z��Dq<F�(