XlxV64EB    2b5d     b10�8prP�eڳ�jG��P"����`��	K$'�s߄�T�ńx�-��@B�d+ٽ\�th#�bV��4���v�e�Z��oW��+��j.�!0F�?lu��,�J�:0�ĔlV&���ڄc�x���L��N{;�ֽ0�Sc�7��.�bK�;��<S�i(�_�2
�@���0c"��׳BVo�����D�o��'&A�L�c��͙�oǸ=<�`� ;*g���q�f.>�H3wa�VW�Z��ta*��<r�(�~j�S��Xo�\"_2I���$�^��2;�ɍh�tN��aȆ�V)S��ɇ��e�hP^�z&E?7�v_m?�q�>���Uv$Q�u$ v���z�ٻ���ؕ�
�+X���P����c�e$�3��x	V� ��n�NH���a#���c�p���؁�2D�1����LTB�Ix�hoe9� H5��CK��3<�gM�'����)6X�N5��o����#w[`�8��z�Xj�������H�jiC�j�pEFߦac�N��anq�Kt���:b�'$����ZtЂ��H'��!���v~��������P�qF����j�_��'e���ؓw�H�X)�m*�$=ۖ�Y$��$
yG�����Y�sE�W���f���_��S���WBI���-(����lߜ*z36#:��5m3U����9s/1���]�����G�g�(��z�M�]$��z���܈��ǡڕ�X����Mn �S�s���f� ����$\Z054�h���T���a�C4�6�p�K�s�k.�|K��!������0�͖��7\b}N]�9���	o��:VNp����@!)��L|�WW�[b�����s��4��c�(�x��$�� ��w������"c[ē�8�6n�p�`�����K�B"HΏƝ�N ����MT�˖�2[���� h<�'������]c��9����j�~���GH빵���tw�����yc���n�V���zaQ���k�����?U��O�.n�o���ax������(�g`�a>,�B,[2�l�����Ø[3���1�m�5�����/�D$��hT��?�3��I���3�3�H^�,��Œ�;	:f
���&�ܴ-/;�_������@��>XH�VQS����~�㿶|�L�1o�&�'A�qd6YX��i���=��]��$y���nOe%�<]N/�=a	{��>�d�F/r��:�� ��耽�C.��t0��R	J1 ��#A�[%�&��+�鱐R��V��7����I@�����ut��_C���	�6��eW��qUP<�űv)}�l�[�;��U�3�q�8�@ ,x����༗`	BO����#���>�Xٙy� ���;Dx��_��G��:��v�nh�3E����*Ѕ.lh����T=/� �i1WWM���ַj\�X�x��s��'����ذ���[�$G�''-=�mxb(2�&��R��&���&�@�/���e�1M��)W���\��4QJ��Y�GG. #"ty�X��mPH��<F��`~4�3�$-n9R�P����׳Q�-�SC[ ,9f���LW�8|V���6>���4/E��{T�8�Ӥ٠�茭���+Y���<k���&J_$(>�)|�|Y-<�Bh+�?5>Ȕ������5�L͔�����F�4��-СՒ�2wR����ۏ��:� �p�<��^��2jL�q��EՒ�"\Gz 1�]�mh�pc,^�.����G�z��1�z�q�g.aS�#1��7���_g����A��+��3Gz���o�Sj}8�_�s�\��#W��ixGca�z	�[=���i§�ى�D�Gv��7���0��U|C������W[E�g�z�T8�,N Q�YM'�L,N��?�O�������$t��ޤ'{&�Y�D���n��u����XLv�M_�FP+z�`F�:A��Bv�f����١X)�V`��g"X�&u>(Ǧ��ۣX�!����o�B<ki���i��s��ܝKO�К�N�n��p?Æ`]3q��wak�
L�HM �6LDZ
匔|� Zg��&�߹(̦��RXk����c}��xk�؁!�1�^���E�
P������6*5ar�-Nj���o,����N���Z���Ɯ�Hj�Vvￋ�����[��͊_e|,Wj�'��;����h�d(��:� x�� �y"W�yڋD�o�k���v�"ˠ��k��,��#�ؘh����ct��R�#\��Ց�m�elm�H4�F~�+�J��à���i�zg�RqCMzi��L&)��:�;���!1�� �K�f���GB��2� ��ϕ�p-ȉ���#ˈ%QyB�Α�X���z�2��|�<r���}P�)�6��Z.m�����ܘ^<_�sBr"\"`-߲�=���K��W9Hi�v���
q��)�^u7rHz+)+�9Vfyy{Bv[CD�K�t|����[�\�^�[Y�!nP; 4a�Q�=	a��B�ro�1�ņ����Ҫ�������r�n�+�v���[MU��ƒX[fK(���(; �D��֓�{.�Q�՟�I�ү�ʙd�a<��S���c���s7�Vl�ZKۼz䀙�����J�b+б��y9$��|1`�8�'��R�E��0��I�-x���A��h�OA}�S3��\�;��B�y�̴#�}����~4Jk�m��.t)���qЙ����7�m�B��fu��
 `L��l�U��7JS�c��J�R�ʒ��[⑆:Q