XlxV64EB    fa00    2850���&U�ȧ�R�xd�=V���}Aӵ��v�-0bwv�#��K��)P�����ɩ.�>��pūo��!�c!�/�yI���xcG��!���c�~d����%���f� s����<4)��7�8�btM�xI;�*�,0�hd@,٧�
����A�+r�����YN�6:u����������Q�hԨ{ӲT(���;6�55Y-AM��
p�ʢ�s�n��L�u���}�dSׇ�<�dB����o�
�[�!�]���Fy�q��(i��δ�,H@� �F��@�h!�]g#W��|�f��;���2�0��� ���u�x"{�]Y�U���y;��<�H�^��QYi�u�{�����`j>�oE�O�'P���,����f#:�l�_&���rx�gZ^� o�����+g�%TSD�욟+F�xlʯ�o�)���Y�5�C������Qf��t�p_��G��#+�o�)�� �'q�3���|o�z�@�H-�$�A�������C�Jq�iJ�,�DR���\�O��4 �G�Z#	C�>Q���mׇ4���;�� ��&��dY��B��dN���`�{��x:�|}�
Td��(m��<�E����x��K#��jz��I/γsl�Ja���xh���h�^o0��#g�mƻ�R x��Ϗ�dh���g�Ify��7XN���ĳK8�4cX�I�����L̳8�'bh��{�/FK��F��~4%�Mg�>΄���[�A0�y^ %��ґ�`��T�NHH�|�m��|N�.�,�w�l�)�g�Z�W�����r��x[�KHt��ނ��
Ii�/V>+ͳ��Hi��|�	��RLw���}!7�MS��c9Mi�mx��m�U����9��2IPbs��Y����u*�(()��<�k(gnQ��s>�ٗ2��Pe�v��Q��"zmZ���T��C%����!�-�gn�IoNuC`���(m5x�C����,�le^ŧ�2S�ےV����Ky}���Ǟٖ�ڵ�20���v`�f�Y|�D[�;����3z!l�� *F����p��l�Ӳ�i&Uy��>��&�ۡN��HکV�F���~�󼰽19���M��v�{��Gz�.���BH��b"�:V�]N�ڄ��1�0����"	���K ���R}Q�<z��KN������݄��8l��1뺌�kO
��L1�<#FO�۲#�L��s������4L�� /R�Qqm$��3���iġ�czƙ���]�[�7H�L3���	r�B�v�w�m)�B��3��i�X�YgϜr��5/xO4��-�d��?NF����~j�S�c���G����/N���Nmo��\�!�ynL<��51�6V;G���ȴ�)lu�a�oj�]:)Ƭ��aO��ad,3���2w��1֕�r��&5��R��bׅnS�EA5ҤK�ޝ#�g�N� ������S�ެ^0��Ȃ����I��>��xp��
ū��J��ϒ�Uh�[y���Ġ\N�3}I�a������5�hO��<�{��b^AV�F�Z�I�.;J�B�Ê��
��ۇ�������_����� �������ǝ�����Ea�Tmb:����
Ά	W�M�H̰IV͙Z��9'{����jŗ�VO|{�қ�0�Lf�e�so&S�u��:�N,��P"�)��G:h�$�y���� �3� ��#}�K�6�	"�O��1'�l�C�t����߲ͅ��m����nA:��;��A�
�_Br���폕���������$��$!�B����l�S�����'4YTY3&�Hu�4P��2�x(��~���lRR�O����*�,D��D
7ry���u���hO��Ŗ����0(h�,�����;���0�D�Z��	��%%�x��;��WV/�)�$��U��nu���� ���w��6I|���B�<Ĺ	=�a�3UP�1x���;أ��23B��ZI��Rp�g5>�"H����y�aHCAzC]�x����|���a�����ͻ���.�Q�z�]��f?�;�ro��b�_cD�V�Ēj��ꕺ��V�Ǔ����f)^�=Mʫ�to�HMn�B:0@�HZb2��h��1���%�9�j�I�SWUpT�-�9�*KpӼ�8e5��V\�a竺�=��N�*�;��ta�S'MN��#%[�.���;�Q�Z�,��������@�,���u#�<�\H�7�aT8�ԃm7�P��x� ����IEĺ ��n��|U;�[���T`#��
��먖�f��{��6�@�ZdP��(�-�� ��晡!��b�7l���8���o���e�Ŭ y���q�?����]�0?KIL[��y��e�;�U.��,���!��5��ۆ
&�����r�/UT�5���úIn���!���{��cF�1!�-Ra�E��v�#<�7x�B����,{uJQ���[�l�|xW�MD�G�g���8���?e�	2�.�A���A��$��$�����H���U������O�M�)�Hv��^�.�u��!� �Pd�6x�zV��2Wq~��}ŧ��?jJVFn_�F��2���
 �ZC��Ȇ����c��$!K_Փc�`����
VU��/��d��Q���V%
�����N�^��d3���e��������}_��g&�Gn����~��I�U���tq�
���&�Ƿ�J�FI����!K�3��ʽ���l�ƃ��W\~����tZ���ɴ�8��;�z�F�����u��ӎ(���V�
���	��mbd����7b��&�d�YR�r�q�@���mI��A0,��q�j�L�sO�R��~�4�����7��q�i
j�ʥ�Q�(�T�Y#p��,38��-V�@GU)�lg��Sl�U�\_6�2vf�IΦ,s��xU�VN!�����TQ�9��e�eW�g�0�.�ǕI� ��]��i�k��޾������a�䟀2���P��.6dq:�F��EX6��\�"���i����y��e�� �`�OI�E���!�?�3���$Y�VG~s�r��KqhԐ0X���f���*��GT�U�������.���J^;���AM��Pu�W��z�G����Kk���h�H����M��b�OYL�*��7Lz��8�"q�����[�����'�r��y
���)� -�[椺w撥�� E��6� ����W+ 1��A���͋ΐ��X,Ng�s+LJG�������Ǟ���[6��-������`�rH��Ԙna��3�����,�<x�	9"�H�/dYLӄs_��Ygd�c�����PZN}*s�K�"[��p����x,��N�l"�.�M��M��F�����v^KE�ȏB�7$H�<��{~������٧��3%��`J��tsmU�����*Ax�X��zѝ�疮��E��uJڠ<k�.D ��k�˝����a��2�,|��8��eNg:=^d��LW�^	4&���y'Һ$%`�PC�&1:���&��M"��DW�W�[� ����,YJ�`f��y{���x�5�d�yJ�攘��c5��\]x�MC�o�Fs�;^$q��1&���\�٣��7qE�#��oH� +n���GL��$��0�`tR�jg�.���1�ρ !|V�����&]�k��I���)��L�^������'E�\�n,��bȁ �}}p��B4}���95|(�(ob9�t7V9M����2:in�7z:�\%�������|_>)Q��l+�V��T2v�����a~�{~��uD1��c���{3}�J�غ��Z�d��haX˔
s3v�85��q��2�'���� ���:���k�O>��g5D�!�i91CF[��)8r�P���H4S��'���*��݌�ev���P�%��wPQ?�|�v�+�5�.�UԴ�-�%W�e�n������������$��8pZ�y����6ŋ5���@©}�ȃ�=��#}�u�7j,$��tQ�-]��^^��ɱ'C����)G�\e�+.Sx�%�%�y�<�8_%�t߮�5���9� q}��5,Cİwލ�Ī� �5V=`0�bQm߈�t��ܛ�d=u7�,4`�.�"�6��jS�X�����N%����N�Na��r<���D^����P�����{�2xֵ���l�M�JVX�.7t@�^�qրU�#����WԼ��X���^m_'��po5������N� ��?�re�R��4�i<�,��ݼ$[��Dmi)�_M6�}D3�8�)���(�]Y�A�/����CEk[��E�K�f�><�� ��"�G�[��y\��ɣj�C�4����I4����[�FaB
$��CG������y?.ܫ����)�� �y���9Y�w�s4��j�шʜ�6�R�����p���07�x��<�0������Z���v!�f}�RF��W���D�@+�f9�&�[\��e��2����)Ü��@���&\(�Z�{��g;�o^���>SI�%��^�ĉp�� D�Q����W�6��U��D�$ �4��.씣���⭣����ԝ��"�=�����uյ;�U�������p��#�(KHmJy,m;*���N�yD&L���!�C����B�0V�\�>F(�c@��]+��p)E�.\��R�	>�b�t
ni4�x(8<zg #l��cm��u1 h�7@P-�w����n�3���
�kYr���.�\�$����������v%�~�[>;MQ%h)��,Mj����	|�$�Ck(J���!'t(�<�׼N���&ӄ %�LX�Kx/��=h��J�����Io��x��H�.	�g[@d�W��k�{t�QO`9�7Nر%�fq3Nŵ��ñ®,�v]#3���&�5K���J�@Y�E������K�,�_8����ɵ"�M�9d��0�/�^s��t���+Z���SJ�[�����k��,�7�+U��Ə��(;���S-�5���)P�d�L��X�"F�9�����S[h:Z��@S�K�F��n]����mv�|e-��`'0��M4dmr�j�����S>��[�E�R�;|��g�)�lsO�8�a �)W�
�D�jg�cU��*zm	.n�������6�>��0�CƦw��υ�U�@������ �e�gw�~="�c+gҼߗ���6<\������j����]Z��� �F�nY��D��͂.��/��g�a:u'H����.B�,c���D3��x��?*��B���RzA�7�}gev��kF�09�-=���n]�V=P�)|�pFk��:�=���6���'�ܥ����d"�Y�&�0�˒~e��������C>ǾI��Qn=A��zL86���i�����HP��1'Xup(��XY�N]�����Sȱ�|[̤����L�k�Wn����Bݲ�������֚�8^�bn�����{ܭK
269��o��Ȳ�1h�ۋF�g/Ԑ%���Z_���������?�e���'����#$�S��f����CO�N��"���{!^�K1X3�),���'����I�&�E��*���zd�Yg�q�S�W��ۆ�>f��
�R�}�=S�,��P�,?o:�XV�-F���Ļs����huU�9��w��U'��]���YYi��.�'�L�n!u�Ö%�#���"��S��p� �Ԟ��N\ly�On��c<��D�=����2ןj�=�x<�\���z	nfb?ݱ�1�S@ Y|=io&���m�ڢ�bVE�L�i��Cc-Ix�_��Ɂ�^*:=���C�>Kи�P�^����l��������IҺZC,�fU�_�C�9�eE��4��\��.��Np��K] b4���ːG ���@����ńq�{4�?�t&#�w�-X>q,�2[&�]P�8��T咷�'Σ�h ��h�;L�p�72�݀RB?d��k]����E�J����C�S;�dk��v}9m��I�f�*J�@l�r�|5�*pHL(��]��nn��q ��-v���Z"J���}N_7$���ߦ�z����~�@<����d|�ɷ(�,2i9w�^��U2�M�AIPL
��Ib
T�D@��툋ܰoO$�$��a���e��� �!��J%NE�-r�0�ͦ;(�R�h7
�@�n�/R��V�H�M�_(ؖ����9�+}y���%ۭ��8e4���+M�g����L�
q�ڊ���.���#|^�)�s�����c�
~T!);���['%�1Z�3����+ߤm�����zȕ�>ޒ��s�;к�x�o��Qm��ɸ��#f�çR��B'!�[�oU��t��!��]�)	y���kF |���l���u\Yc�Da�~���=͉�w�Bd���<pr ��*�>Z�\�[�q\���H	����i�=Z���FߗQD�W�o�l)����`�&�T��.ҹ��j�Ht��OO�����4��@(��ĩ�f�/Ez�ur�Z����Ia��e=��Le�0�W��
�Nk2t����yR�"�Ti^��4�l	&���	����䥯��Y�8�%��f�K���`K��ͺ�j8��L@!�����(1M�D\!G�����6`�㉾�_��.���pY�w(�r�I��S"�-^�'�!��־h��|�{���@kqc)�48�n��G-�'Q�y�̼�3qg����Z.\^Awd�ď+!i�^�ة���?6�����B?��d5d&���h˞*jG�޳}�&�#��^�UC�����unΰX��J4�T��lՙUBOV�i[mY�.���A�&L��4u:��z5䝗�����J�V��v����s\�.b��d�rɗ9n�vIѠ����m���� !K�GR�=��#�-�a<���z���@5�D����*6O�&tڎ��]8GZg6�������xPY��"��5Jj�� <[�d};�몀�� *~�24�B��Ӈ,�>u�T���n?�0��F�㼥y�Zn�;W@1׿���ŕ5A=$�^�<���2�C���G�~�S t;;��(����ړ�.W���4R�qH�������Sq3�U��dq=���2��0��DF����Jz�������%�2�@%���'�^�.�՗wM���\wٟ�#�pҟ�����"Lu��@Y�!��U�e�A�5�bʒ�fL6�@�����n3��O�"�А�ݎ|Q5I�G�H�n�DXek�v�r}$`���h��Լ�1�����8T�����KݑƱ �
e�y�� x������M)�������{s*�߶�7I��w�#�)�ԁݕ����K�l���x%���	���0��!`{�c,��g��P�5z$8����������
T���Њ؃��ߵ���]C5"�y�^)����}����ϵ�X�M���|��-�!�]���a�Y]�\��������,a�+��sX�㠔/��{o������;�4ڼ����Hj�d�U*(7y�7��vR}A=@���K5�3�+
�A��U�Ӈ� 	Zk���CfN�Q������%��:�]҇�b�x��gp�.K���ȉ��a��m�r�B�߁qϷ�}
���44D���:݇\	��޳e��O�,37"���l:X��Ev�ʂ����8��BuG�w>*�ٞ�����0@l����݉T��KB��H��t�oӹP��ɭƖ�ԩ�>�ۜ�,ҕu:��0胱��jI[�z�_�����c����;�(�B4���w- ����/p3z��G�<�!0��n�?��3�HS�]��.���
:3 �6��D�M�UyԻ�vB��U�(}�9���[�����Zk�l��J��w7٥���A�<d��q�d���2��H���Z//�"���%�|0�/�6�Oz=J��pj��@"Փ����9�]U�`f�����$���=��=�L9RU���[%Dѓ�KL�Kos�n��_�e����t�q��a��U�\�(�'�j$%��`M%.�XF�]�v��6T-#Cw��ߨߦ\?���
��
P,MZ���;��n�if�;�3��Uհc[���fޅ�TB:��񋎾#�4N^�8���e����B�jhSPs�*r��
��}�mA���Cu�����K��j?���Irل�@p1��x�'��1
� I�4Zb����C����t���})��<KcU�7+�_43���!�w�k���s��6������0�ڀB�ꃑn8h�W��,����h_���-�T��5�U��L�6��ڕ��5LY��Jk���<vy�t����#M��������D"3h����I_��|�bM�$)���� ��(���c�7�p�4mX��蠴/g��uy��f]7U���D�ďԎC��R�N�w&3��^�_���]^rfxM��;��]�/u�O|.��������f�.����%8+d;�Vئr���p�2Zr������{���^6���'�~�e�C$����"58��&��ȏ@s�\���������1>�c�\�ؿ��� �Te���IV_�hIb��v�����'�.0���S0��M�#�}p�Hi0�P�b�66L÷��9PV�7�Z.&܅�Ѳ!��u5�`C�=��o�6� *V���/am+���(�b�G(߹\�g�M�<�6�
hPG]v?��CW�%&'xf��9���5�v "���`$8����[�VN��	��Z�"���~qx�]~}d4{u����e�?ݷ��E zW�7� ��,Ѡ�9����E]]&f������^+@+χ�J�t���U�|RzW�->�y�/�q$�k$�<u&^�6
� أ�V+�e�M@?��p�10Y{��)ugv`\��>i�� ��A�~d}�a�ܝ[v[����0��iL����D}N�	 R %�����j��=��h7W3K�m.���� ����+J��NTONҳ��-�B�%�-fnE�e�-���@t֔�^���0��o�t��2%=��n{ҵsO(�	bV�z�7Z�`�&m�,�	@E������kS���EL��ϸ���c[�Ӷ(�B.��\z�,jm��h�I�G)�w��{Yq�?
i҇q���J����eA��
�h�uS�Z͚���,	1��� �!�� Q�Q(P����C; �d�@.�&�FEY�54K��P ��칼S�K�H�/^֝W�f�$�FLz�L�M��!��k4��H��Tm�8w�� B�֩��g"�=���F�$y�fT"<��и�+�AZ�>3I��XOR"�j�v�H���$��Q���\;[���b��ur��[�/��<�m������I�)�"
�y=�;��<8f���A�?��C������?\|�Y��w�1����E�-�s&Gl��|'�.�JyG�ZC�����Yx���K&S@7����*u��X�T���������qLn�&�aC[q��'4i"?�H���ű��9EN���A����ҏƸ����[����'F*և��B���nvbƭw�ߘ�-�dil+)�fw2O��t�t2���M|)2�0�`��z�|t������q�'+)��#ߞ�<�5ک,�Ѳ\��FzJ��F���<7Ci�h%k�z�S�hk�ElۿD.^5��j���C�<�*�l���A���]����-��B���Hu�;�$��1r���_��q�v�z`ЬB�D`i�Ϥ���Fn	/B{�MX�L9F2�q�YMc�3����Y���82-�U�E��������f�E�#$1��i2����z�
�g���'#[6�=��I�"�~�P9d4}��*��� � ���\��O�K�by�i))2���)��*1~�o�N�B�|&]Ĭ�"���s�0HFہ0���V���&j`�QȎf*�s�鷽�vf.����xYpsX{����__T�Y�ls�t��&f��z#� �	,2j���*�~�zؘ�-�*|��N�)�RgmӦ�4�~k�4=rz�y��v� ̽�$qG�(Jmx"�$S��/F� [ٳ��>xs:�?i���b%<e�� ��g`��dP�&!���.�|�	�re�
 ��?0^�B�ڊ9͈�v˪�@�6�ё$��~����kf�JuncR�%��$l�ۆ�9LvZS��O�A������
b,
�t[����~z����H�E-�\�o�"XlxV64EB    6c4c    1450#
����)�o�X�J�7�a�2Y�]e�6��?y&�{�٢vn����%N����)�;����P@"�J>��ڝ�MU\�J4��!A�QK$�]�7�IM���d�-l=x�_F��-e�� r{�Gɛ�&��X~���x�Y���!�"ڜ�?vs>��W�c��R��q[|�|�p.Qx�����V�Z���pR~x=x�\������S�W����H v���^��U�g�_O��]�����t`G�����{nI#A��: (�'�O��j~����!Yz�vg#���x~�$(��W����h>P]N	�<kH<��J��� 5s������/�{��(��g��ծ�*{��۶\Hb@��՟ɔ9
��gX,KV$�7E�남.	F���0£���S���:f������S'���/>#C��FJP�5)�N�
Z��d�P�����%W����,�ܹ�P�����h�}�Oգ���:ʘ
f@ŗ�Q�*��[8R�J>/֐w�)f�FQJ��~��F�4b�󊩊ϥ�U��"A�؈�	�Ub�WK�E�1�x�a��M�"*��l+�6�`^��*���4�#�8��[MB��8�5Bqt�,#�ZF�;dX�ʝJ	�U����� ����Ānk���K�~�n��}e, ���V�{��]����&��L��E�j?>�cH ����M����V\>ۨ�O�lE=�yg0F��!�m�e�b�ӿʸl��aE��n��P����S�*��D\�`�8p�,�ξ�}e�Jͬ}0%�]��!�aK�����sD?$k7/t��n��w�Z�Uj !gh]Qƍ2��FJ7�w��22'�8�2���#p&�+%����v%H����\�0�:/��[u���<�Y��-UG��`�c-Dְ���G��������D�%��8����L��v��V�	(e����@�Āp�إ��^J�5���d����q="e�H���R�,�HB~��&X�F�C�tU<��'t��w��8{�M!V��U�m��`�����es�<N>>a�&p��n�^���T.�ծ�أ�%���<?ԛ�"��fz&�����{��m+��ʟ`S1�-�x6"ܓwΖl�"w۶f��j��敘bȄ�C���CiK����%���V��J��`֙�XM!�t^����=�5M�_w�g�8=\RG�YN�5>趏���ݴ��	,�����Nf �M�A�<��B�)Gt�ju��4^�̜�]�g1�9n몁z��/�̣�_��R��e3���-<��Ź�,?�9|L�j���&�`d1�<�u��؟)�I��Nʎ��_f�XA?�|�-ي��v�1ߑ�B�4D�S��<-����,V��@b�h�r6_�5e،;jT,��*XO�xʋD�*m�/QP�@���d�Ƥ߹�	+��e�ފ(ZkW鯹d}C��=}�����W����i�|�E�|ӚW�V�3R�c�c��]�9-;)2��@AqTFk����MS;��-,vbg��� X"7��B�����Js��"5���z3BB�ks���88�%�L���t�
���^����L�A�s[{x�n{I{�� ������Y:�&7��d��o_�L
�[�Sw"��Or
������L��0�IT�V%�U���j}([�ҬM�>�(�\r�� dÛ$|Ŗ=6㍰w�MV.����AA��Э�MT��5[l<��3��F��@q����������7Vk���d���xM~�!���t9$�6,��>�8�ސM�jO��qO�� �?��s>� �_/���ЮW�Y�y���ї�\��[��1y���"�V�u�b����v���.�+�Yv�{ߞ��
�) 5�����Ck"ݭv�_�.L����0"w�%�Ԫ2�̴3􅞭�^���,�{���>ҡ,�	�!��������a��=���v����nSOKUح�u�1��g����b}�i6]�)�FX�*�22�y�5�71�J����W����	�Z��J�{z�⅁W����}�;�]p�ى�?�
H���z[~?�����\F������Q)����Z6�jC�����B4}r�2eܳ[K�UZ�XJ�z<�����H���U����B_��G��~�E<Sya�JCX5�a�b��r��
�_��/3ϩQ�+6���O�������R�`bƷqJ�I8����i�?�!T�(h��B�e�6I�T0���e�F�]��0�io���$���,4h�ɏ6�d����ݰ�P��ҘBg?�V><�,��J����rµ���4<P��Mk6��m�t������rdyE�S��6׉L*8�1(�N���*�_�9���3�W(4��v�`7���)o4c��Մlh�T7��ܲ�M��䒇�k��R^}�Z,�$���M�d��ǆ�$΋�<�ݝ��YeI�:�n��R؁p��i鈁&�zS�ڙ2V�}<#��7������)iȍ}j�(q\��,�Dp���7`�!�9�֒��yn���jO�! p�v�6�T)�*M˓E<�	�y�bzbr������۴GM�N@�p����#��6�<}PԵ����2خ���Oe�H�=Ӏ��:���{��'��1yʯ�:���vk[{�P ��^��s�a1A�Іfԋ���������)I?�\��G�Q���L{���r$__U����h�R<ֲ52��ca�����p'����&�w��-ED�/�	��;hC�QҶ7��{��|l�T[�=��
m��1�0��H��Vmq>��,�͹�u2�3eo����.�#~��E�5�!E9
�a�|��3F���wXדr
�2T$��a����k����yh:�1��1��
��2W���Q���k��34X+�xbt���j��Ƌ�5�V�>F�#��
~��y���� 4[a�FAh�����J�_��.YMr#��Vjq@�b9�\e����,���a�=��9-��D�Q��|����v�ir�)%�vlB��f�����%��v>�f���7i�i����E� �|�R�L��(8_�R�-��I+-v,�1�/��-6$�����@/�'�ma&�ï*�]�n�o�j�*-��l�M�F�$O��#�C�Nv���=��Ji��Y��IX�{��e~��z`Vy!���B�{E����DM0³\���o�͓:m,	Əc�=�{}���!bVː��6Jj�}��z�H��3��Osېm
����ڬ7�?'ɀ"%�m�f��	!��ң�G�����_	�,�e�nlC�4J��VC7r�Y	ϿS�y@<��{��<��b�EF�^�R���e��u��!�@�]�i�r�EɈ���4�c�E��)�/a�R��w�V8{`�W�@��[�j�Ӎ�x���˼g�� ,�|PD�^��P/�￀I�H�|w|k:�Iw�?�AT����@�]v���UW�5Bٜ'�ϭ��?ةG+����;v�^�	J��YvY�h�A�≯�ni�����kK��IQ�i+ [�`�P;#�F�01�}�1��\�����xz�.,����^m�)Z�1j���%S�[�tM����룬�8o"�7� �ä�v�"l V�Lyc��ax�aI���
|�*=[6��)]�����g���rFt��V#��~����ȳ+x���˯Cf�Dk�y{��EI [ � L�)M/�����c\"E�vF��x$�'#�Ѥ8���K�V��`�����"��F}@٧�R�{Y�zo1��0%��2�Wɐ��q�Yn���wM���z����_��3u�XU}"y�a�<wyqسZ�HW�7 ��r'�_�0������U<�jQ��;��͵V�g;��&v��X�U(�em�+NV}y�&"�pI[w��&yz2-�~eE����8$~1�_��fb�Ҕ�C���i5��P��3	y/�u�"^�',�(���'�g)�#}��}���P�6������W
|��Ճ�5��諄�*�_�����ޞU���Xu"��G3�����->�'=��|��l#SG`HjBc�J:
nE)��|��Q��v���Y� .���3�ne&EÇ��[:W�CW_P�S�B|�ٖTv�Ju{AƌY͑���nZ_g�ˊ�U�a���q�|�MM9�$���^:gR�J�����j�^I(Ӡ�?�qx�h��r�^F��5�_7Ð5l���t�u0)[���QX-�Id��U��*lJ�0$X<�@a�=���+2�;N�:��^p'*�.]F�!!๚���E�"����J���\�?������98���"ۘ�.OAu���ia�.���?hxδ���q"�J3#L{Y�RE�����Jʓ�ñu��WT^j�O�����y"�04#�w���?��M��T���=�,]�i�E-�.��.��-e�P�1����E�Ș �^C��ܝ��~[O�}sK=@W����L=p�9��^���U���*��5W�nf�E�Ԧ�`�d�
����x"O��>��yQ�w�sb��C���Լ�	͘x��"�b���8�R��A�<�L�� K�g�X(���y4�ܰqY�� m2�;[�\��ݞ�ތ̹��)�gpu���\��<TƯo˓�������D?M_c*��0��������@�d��Хa�%+�z[W��Z/��a:�K�N7�ܨDF���H�_ur8��~�/��̬Z��7DȒ����I;Әe�w��$�ޒ�ҷ4�~oH䅧m�{1(�2�zʩe0g�^ M�ı=�83�!F׉��?u�]�a�U�h� ',�a���p\%Z�l#+��z���X|��Բ	������:,�*n���>�U\��T���T�"\����z���r�G��2�M�聻R�:�
�Ar,�ƶN�<��T(�r���7(�p`���1���rPQ�d��@�d˼�/�}�|����T���{�����K�� 5rF�GGl����N~���~��$�����z�C�+ҹ�$�fE2���S+\wk�>۸�N�r+W��G�����l��w~�YB�Zx�Tǭ!��C�7����Q3�g� A��+�'�pm�����;6�;H���z�)