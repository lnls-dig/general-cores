XlxV64EB    480f    10d0Ǎ���JZ^w+Q��x�L�!�@OKD���A���N	�Fn?��8Π�6/�}��+`�X�y!�*��L6�����Kw|$��Y�;$!�cϑ�YY��K�d-U���꫈�����Y���)��/b���V�{�-��� �2���R��VJ}���ax���a�v��!�p	�0��\�t�2w'�@�n����Ύ��Z��kH�5���g���k�F�b�Q�� \�ej�����T���Q�v�v��T�O��PucV%&1�o���H��fs�1o�zπ{�� ��oເ��*Pj�1��=G��4�����`�
-`C��	n�ͭ�����:�͌��bQA�a�Q��ٕ,
� �Sk�?� <�����.�5V�՝]h��M>��oJMn�?9��~�]�������X&�����+w*/ ��G�_�$�&I����|�L0�4'hI�4<#��kM}:�$>eBM��;�ϱ_1�fј�d��o�{��Ҵ�F�2��ʓ
��\�4 
���ߥ,�~g�_c����8g%BY:�F��E� �]����U�Ȭ��#�.���_=�Ӏ�b��9��T�rb:��`T��Jt��ڋ~@�q��^�P�$/��7
�L���J!��;Q���^����&l��(���s����Rc�,[>�����+��  ���Wʠ�Rb@� n����Qc�5p���О�0ta�Ƅ��=&"9�W&D��؅MD���,�a�_�n�9��C�b�3�9>�sR~}4�����/!�6O�yY�0�n&�	�^Q�&�p
1����?t��r�>�Ö���h��?+ �ˍbR	z�Z��χzD����J ��.^/�����[j�˔��m��Dp���rL5�����Dَ�n<���~혖 ��5��b�����MS�0�c�`h���%�$g�I��uG�3a	C�5�р�f�Xƈ ��DYDKN��e�Rȳ���$���*|����Ȫ�aQq���1�<5�O,�v�t�@�碲jbs�Ğ��c7ɺ�n<��*��}O� �:S�I��&�D%��G� �#F���!*�E^7����"�f�X��=G���iX
M��ZxÃR�T��ntq	���X�j��|�)$W�����'Kv��w�d����y\8�P��Cm)�6�OB���*��[˨��~s�(��U{Q�#����˅9���И��/ D�o�oZc};8	����������v	u�d�m�ݣf_,N!�<����`a2�C���'�t�O�@��^;�΁W-�*��5��q��}9���XUS��G���q���u�/J�M3yG,��S^G� �s�����@�7�a(�5�x�.z?:����������t�œV�ع���O�����=���+�A�\"A�-�ׅ>OL���ģE���x*q�o��=s�giI����~)>���1@�Z�Ѫ�7�qw�^P�ո�a�O/�OCP���;G::)kV�Q�'�b3�[�Ыuz���B�1��0�"�JT�t����I�e��E��;U>����#	9Ɵ�Q�&z��C�J��DB�!DV�Od��{�Ve~W�7�w�ٸp�Oi9p��<W��ݺ���v���MvTzG:���k�O]i�#Z[E4�kP�7�P+�4�,�&���J����XՋ���K׈�.��ӌR����1,~~���0joح	�̠�bQ`Hk[� �c<DDV��NF�]V:c�`�)d�gA�hD�²���^ �'����'��C"}�h�	A�����3�׾������S��j��&�P;�C�1�7l̗Au���ͽ���ʺ���)��N��;+���s[ �x�"��3�}��+C�|b�}��D�����B231���a<E�BR	��joYx<�Th<��dY��> �O�9i(.[CClM+��R����3����+o�Cf���5;�7�,~T�Sz�ۣ��z3��P9F�L���zY�y"�p:W�$��z?�R�9���i�&#�*{
�^�_n����dw�U��G��:75V�JT�Ct�����	_�|~�T�v_[��[�G� _\ARo�n��XS��-fs-�]v������j���00і;�d����O�kV%�0�
�>i���Z;���s���MÊ+y�ϝ�}�׏�w��N���ɥ�zpeA��t�1bҎs��vu$���/���c*_|"w)�hsyf�Q��OƂ��iL��6S������ӓ� ��8[�:q�r#�LFy�m�fS������̙�,�4��@�G�#bv�2v NozE�����Ÿ
.�/��̖�1/��5ۦm���L���m�|h?<O>w���an2��IA���x��C�~�4�u���m.�T��F�H�)#w�l���[��(�Sh#�R!��yOd�g�I؝̪��� o�0���aH2q_M^G�����\:��K�E	mP�����X:j�w��~
H��=?��{5?-�I��K-��Rg�мr�B߅<�(����4�$�:�~�����Q���:	�&�낺�nE~tV�MH�&E0䉸��i��&�s�JT�ٛPa>�Y���/��g�(���B�l^4��g�VU��3��&��QAcI��?������񛣥z�F��L��l�Y,�Ӈg`W�TG��ؕ��gwv*�[���8���浍QE|�ptn�����r�8�~uL���W7�K��"N�ac� ���<f��];,��m���F�im��U�æ�X.N?Ik�O�@2���X�:�U��8�J����U��;n�g{�O��ӡ�C�YdJ�g�E<�l�J�hR5bJ]��9�ҌQ��zO�!k��bo�)U�qb`��V����#���J٥W��m�*�g�o��N��K	� 46�/��>3���q<%�A҅/xc��`h=�d؂���κTP�4���G�^���>��.������5X��	tʊQa�@Rx�=�>q����{Bq���%��
g��T��H���T��&B.�J�?0=��D��u��z�HǼ�t��(W����k+Xx���?zN��%�E_�p�:#Z&��2�OsE2��}5n}�	O�3�#H�7 ]�'6�R�H��0|b'���%>�9��T]c�Y���}|�t=W�¸�6u�O@8y��Hv�Ybz��oz�����k)��y"�F�����Q�/.��)�қ��Uߍ���b���8$�y<�,[�4w�E2v�`����R���ùQ�b?I@8M��ZV�`a��]��g�9Fڭ�L�GP��d.
����3na T��K7�=W&��(�h>|��;��h�A��%V�,�}�qW �'������Jd�F��r�J#������u�17��S�2θ�cO�C�+b���7I��y+��������w�y(	��VH@?Q��E��P��[uM::���w)��l�b���L)�P������q����\�7��}�V��DRMu��?`u��Xnʵ6��V�*���2g�����-0!�Qo%Qc�-���Q���d��]Q��NDT�;$!�4����2�:R�ܻ����w\�8XD��𲫟��L�wԒu��.l1����P����M��BM�/��C�P��fOf��?ϝ�n3ѧ5�B����¦�Z8��e�ܕ�Of1�Ɖ#���57�9m�}��s6Н�������`�G,��c�n �Ic�1�9���s���8z�7�m��9A���]��xz��?�<����N�L�?�t�����9�n��N�KI�eޞr9��E�B��ʃ^w�Ð@?�G=�<l��
��ؼ�4� k�R�����Vة�	I55�=�W�k���ׂ����]�\T��ڦ�C�F�B	붨�
�v�*�2��#G+�4���F"�8���gkQ@h]����2ǆ0e����
�{w��SC�����F#��Oz��F���\�
���?E��C
�}M�'�ٔ2��J�H�y�
�pD��xYꉮ�C\����V���)cH�e����/u �q�N��6�����ß"�wn#�C��ӣ���.R�oi-v���7���]:G_�E=��r0k*2��늪=P
���+���QS������F�rp\��P�LU㫯7��:�ӧ#AY�ǧ�2&s)
�s$��]���v�!1��`�K8f�<�d��b���0�j�YU�ӵ� N]�)��w2��ûe,�H���"5��oeh��7�.�/z`�