XlxV64EB    5366    10a0�'�:4�3!�=g��{!��5D���k��+#:�ML���������Xv�(�ż����dAn{�;C �~;���&</\y�2�oS_�.�����K)G�5R$�&�o�"����<����<���d:g뎁O�1�g����+�󊍿<%�����G�d*R�� �Dd�x\�V�ʖ-�EQ�;z`<���!8`�3���9�l�pҺ��R�E�'i!H���v��@�\-	i�i�&���a�����}#������/���6���3F�}�z�B����,"+e�����5�Fx$H��s#`3�>�n���l<q�l�.j�e��ѸS���n7q$],+��`،Ђ7#����e�>�*FsD�/�ʽ6�L��c鱳gg�Ѻ�}��>���"l`���� �M�ޖ��� D�]A��O�@��F��>u�&�Lciho.�T�<�`['ɯ-S=&qB���e�B%>fQB�{�Aii���RL���fr��)�]���|��g&7���3;�2u��$ʱ}�ʈ6d��=S���y�hr�q�?�b ���yu�ܖw����@�9�#4���ُVGLN�C��î��`��Fg�#��e����'�9C��5펚l̩��}z&w����4�;��i�����Aq��-�0�#�����޺�2,���O�׮��e�S�u=�Q���f���[n��,��q���9_8MU���q�p7ȃF�u�̏ML����#��\=EbȹR��u�0%��,g7�ji#j�HU��;v�e���s�tc<S��P�u�����X�gS�\���?�z$���ye��<]��
��xR���K�}G�n��*��olh�p3���	��$�I�+�W�I��6���$��B��py��i&0���(��Sb(�m�I=�:!���v������Q{�� ��~v_�0e��G['	����`�������7c��VB�������D��Xv�~ELs<>bH\���Ӱ.�L��Jۮ�@��8`H��A��4��W�:Kq��v��������MB��T�ˉ�I�O��d�q�j��k�ZL�.=�|uŪ٭-�x]�E7�/�5*�Ѹ���PB�����{tvg�m?%yV��X������Tަ/"�3�V~�k�+��2�k��NX�b�^g.C.r\� ���u�=l�]�8i���D�ͮ\����8��.wg���[p1 #��Cr��D+�����Z��0�5��K1[��Ǉ��F�$Ɩ7ASe��U��r���Ȅ_��Epz�$�`��=E���d����쥩͏At�ת�(}��~�q�=I>�0=0�8�Y[��,���e����$�X����S��\�&p'�	1_����E�Ū>��=��r5���}B*��<�ޚ�K�/͇aI���g<��r_%<�8��We�o�1���^G��-�¥����M������Od���jd+�:��ʜ�3��4JϮ�\=Rd6��aA ,2��wɚ��k��'�M_�'��:�Qu�t���J"hz���H����E��m�?3{�s��i2�)_��^ώ���-��������|\��d���f8���ڨ�����D�ߍm��z� ����Tb���CB�� �l"LV*$�o��b�OØ�k\�V�PK�8ʻ���(��v��d���g���W�Ðx�Fh�L�cZr&����B�Ŧ�\T��0lHB#�o5��m�E��}n�j�ǧ�'V�䲖󥐷��o���%v|�R,3���c��^3���r�.��_j���sJܝ����ڒAm�DFLN'_��	8m?�Ӱ*� ��+>~?:}�[�̜HH�5h�ڷ���F*�� (3f}���
8���佀��:hG�$ʙ`�M1U��O��%�`Ո����R� H����ɴd7�����l*��C�8�<���r��0\�S�����i�ȅ��+�=����q�u�AE���I�ZW���y��W���"!t{��o��zN3��5�0��A�	�*�E�Yr!�E{�j��B�V�A�,A�.��E�_0��^k�uˉ	��f�L1k�)A�=��4C=��U�.Qh��<�,��Қ�fky`Q�=7��?+E��Γ6�L0Z%�8�Dc�3W���#S���tPC������		��n�9�P��=įqv���T�)�����ӿFͩ��:�.0�b#�Q�lj�Q���ːP#T�r�!���;��B�M��A�b����q��Q�7\����+  ��ܣ<�9�*��#��'�D�n��xzq�q����c���W�3E��r�_<S-Rh�N��OW]~�.''��FHIm�|��w��*���-���:��잣�4ʢ�AG*�Qy%G�6�DW�i-ѝ!��;@I�y�c�7�@���撡Z��("���r�rl.�uYHH��vR ���/��C
��;������c�0��;2�&��Z٦,l��<���������w��=ߤp���p��?kl-�.-�if�7��1�S��yԬ�7.3�0N������ҥh&�1ǰ
�i��؉Q��&[�p�1FT1������#Y�цbf�T�0�z��5�?l��f-�V
���3�}�Ĳhǭ�B�G����{&��VN���w���O2BY%��g�˽���*8G%�ֻj����0@�\�,���#E�xF{��7��.�ŵG��%��+��N��=4R�]��p2T/A�q&�.��g�vR/�h�_xɹAs^�|Щ�%Mb��C�×4� ��ha+��L��5x;���Z�¿�s�أ�ۇ3^�ԙA4��ws��&"����c�y+�Oͥ{�Rg*��&�]"����A�����g_��9%�V1���i���f���?���Sr��'����z�7�@�Vi$��5N��W�06�sf�Jϴ�Q��S���h�����!�H��7��E:�şGy��ȹ{;�چ]���>hJO�����\�%2���!�UPjv��֍��?ʰ�?�t�@��4�������'���2��+�-��W.ݘr�<Pa�Zy�6Hȟ����>� hZ�&/ⶌkr��U�^�����k9���P�O����d��O�d�2[���K\�F;��ƑN��n}d�/	TN>��%�i���ճ���n����C�\q�y)�mv�����:O}�Y{v˼N�b� �ы���>4P�P	@P�NjT��oQ�d�|���(�_�E�o�0�R�!V]j��Ӻ��3#������IQ=fD�TH^@���X̌��F��a:`tA������FQ�?���SW��
��PV(��/V)��_�zi<~�f=D̢��8/�H�����L*�	���P�a ��ʹ�z�q��/��S�ˈ�����Ǔur�1_�X��fs���x3S�9��Vy�Ǿj�n{Z��~'�$G�Uc��ю����[�
�X{������4�����Ez��-�ޚ���ٲF֗��D��z �'a8��p�^�fHRj�j�?�� )C-h�]Pk��$)���&�6��1gG�^f� M�$0P5�����6�$�S0\0�M����V���N���I�"�xF�
���P��7��!_�U�.��Vk�pE�S_����
9-���cqԏs�ߙ�T�Ík/��e'�UQ+(�&6�u��ܺJ�����-�&�߅�c���iz��n����+�3�گ����^�@�2�|����vN��I)�iDRo�҉u2��-�(:y���7O1�p�Hr6���(�kT�8jtNt��6���X��"/�[6q�I��T&�
�۸�5��sP��ϸ�T" �n_�Bܨ�vS�"TYX�q�F���N������J�-���%ܼ+�eCf9�(x�Ds���)*���/C��y��v�.����%�6��r�e۞1P�5��˸�[�q*�O�����/���NF��笃Rz<-���vU��1a\�[����˺�4�&8��G;�`��Qrh��Ξ��9EYn�Z�/��L�T����Y�v�V�'C%�b�%�
�*������W�U�'��d"���Wab�~y���H�a�$-x�8�=��E�`��wb��;���)1��(��3M��O��A%�}�.�v��S�_��Jj�Q��}:�>��|#����D=I���G���&�������