`define ADDR_UART_SR                   5'h0
`define UART_SR_TX_BUSY_OFFSET 0
`define UART_SR_TX_BUSY 32'h00000001
`define UART_SR_RX_RDY_OFFSET 1
`define UART_SR_RX_RDY 32'h00000002
`define UART_SR_RX_FIFO_SUPPORTED_OFFSET 2
`define UART_SR_RX_FIFO_SUPPORTED 32'h00000004
`define UART_SR_TX_FIFO_SUPPORTED_OFFSET 3
`define UART_SR_TX_FIFO_SUPPORTED 32'h00000008
`define UART_SR_RX_FIFO_VALID_OFFSET 4
`define UART_SR_RX_FIFO_VALID 32'h00000010
`define UART_SR_TX_FIFO_EMPTY_OFFSET 5
`define UART_SR_TX_FIFO_EMPTY 32'h00000020
`define UART_SR_TX_FIFO_FULL_OFFSET 6
`define UART_SR_TX_FIFO_FULL 32'h00000040
`define UART_SR_RX_FIFO_OVERFLOW_OFFSET 7
`define UART_SR_RX_FIFO_OVERFLOW 32'h00000080
`define UART_SR_RX_FIFO_BYTES_OFFSET 8
`define UART_SR_RX_FIFO_BYTES 32'h00ffff00
`define ADDR_UART_BCR                  5'h4
`define ADDR_UART_TDR                  5'h8
`define UART_TDR_TX_DATA_OFFSET 0
`define UART_TDR_TX_DATA 32'h000000ff
`define ADDR_UART_RDR                  5'hc
`define UART_RDR_RX_DATA_OFFSET 0
`define UART_RDR_RX_DATA 32'h000000ff
`define ADDR_UART_HOST_TDR             5'h10
`define UART_HOST_TDR_DATA_OFFSET 0
`define UART_HOST_TDR_DATA 32'h000000ff
`define UART_HOST_TDR_RDY_OFFSET 8
`define UART_HOST_TDR_RDY 32'h00000100
`define ADDR_UART_HOST_RDR             5'h14
`define UART_HOST_RDR_DATA_OFFSET 0
`define UART_HOST_RDR_DATA 32'h000000ff
`define UART_HOST_RDR_RDY_OFFSET 8
`define UART_HOST_RDR_RDY 32'h00000100
`define UART_HOST_RDR_COUNT_OFFSET 9
`define UART_HOST_RDR_COUNT 32'h01fffe00
`define ADDR_UART_CR                   5'h18
`define UART_CR_RX_FIFO_PURGE_OFFSET 0
`define UART_CR_RX_FIFO_PURGE 32'h00000001
`define UART_CR_TX_FIFO_PURGE_OFFSET 1
`define UART_CR_TX_FIFO_PURGE 32'h00000002
