XlxV64EB    4349     e50@�������e�9f0f���?�����u����E0�Q>ߐ "�<���\��q��V�k;���Ղ��+&n)�@e^��G�E�nR�eJ��U�&WW�"��籟�Q	����K@�N�O��B)�,٬��HeWbm��t�:X"����C��{R,�d�hc+�z"v}�o$�A�u��!���В�9O�������Y�FAk`H�|�$�'��#��x�g|��L��D��?��ԜM��X��d`E���ѕ ��MRy�X唇j�$D��LB��y���<��?��8��E���!V�H�k%�f�����N-���0
���*nk�`�I�+�]]�2[�f-��Bb�"a���'Gp��=>��o���^�K�T��UM_k�����5ބUN��F4!1҈ۘ�S����|c�~'��������B[=΋��L۵eA� ����Ǵ������%�"�>�����j����dp�?\"��i��bi��ʙ��Z�G�
�����;*���@�N��l�|m�E���v��f��1�F%{=�� F�˜ �4�x�_�fe`+vjK3X$�Rfl�P�`��RjSo��7�i����WN,*�(a���zS�g֢2� �0Nq�*�H�5f.�Wo+n2����ᔪ�/U����v�M=X�(5�N�m��J��K�t:��-@Y���_����Wp���e� ��=!�ab.����w��^��h��1�����b��+�6�4�O�^3�ͬ��� ��ڋ*E�m��<Eٮ�a�~6l��Ni�HL|)5Ŭ�r���_�}�`�y��+���*�S}��?���������y>{'�Ar�'���\jL���d�
�!�9����.�>�h ���9��]RM�TF"���=v�sܔ5��Q�fYX61"�>8q9�K��uX��f__�^X�V�Y�|��}Ǳ?vr�����c	��~��kX)�rO�"V'w��O1�������%��&T}�l��x��e�t�|�aK����K������YX�y����2��]|�D�����RJF� t��~\办G$v�l�$����cb�(闝q�y��An���g,�Ψ2��$�s^�&rȄ$m�vG1�j$��@�~z�?9Ю9��'L1��9+C��{�j��,ZN0An�����?mR���Ғ ��;j�P���;�^��~���Y
��Z���PT���$[#6���5��-�ؕ�F�K��5�ؗ�9��H8]���wVȱ�3-ɧ�FOtc{��$"*&���`��0.$�3^�Ll0��"��:%x]૝��^�@��̷���X5{�D ���<�&���60�R�N3���T��p�(1&�
�~�!x��ߟ���P1�Rf�m�_���0G}Ѿ�#i��k����#J�����Q�c�@9!��Ѱ�f>�Vݎ&��+G�leF�g�7T\�(`�B*2�վ>4��#�1<��s��3��hSJ���r1�J�O���.�t:��5�M�3R����t��d�� �� ����}��e��Ub�o�Lͽc��Ƣ�4Axֶ��f ��!x��6����l^>�Uͪ�͠��8ԐW���ϡ��-6���"=�=�������^pk���鮌���W5^�V�=�F��!#�am9�܀�f:#O���������Q��Zʞ8����~��l6��4��Iv侽P����.O:#.�xL���J�N�B'{:���1K�' �u�IQ5��u)�F=b�@Ų��\K�zq�}�fލdsD����Az��"��S��ٖ_7.�Bz��O]���������R���u&^�S�2G��"k���Vw��4�Q�xꨱؖ I)oc�HĚ�UG°^]�!�#��</�͙HC���,�n;M�-���U��\`MBo�Q2S���և`=����2�����9>�Z���yǕ�b�tA,�\o���ؠ�Ō�i��rY U=h �����Ĩ1��!�Zy�/Z4�Qx��]��+�U�����aCw�I�䌧:͉ �k��Z�Qx�+��G�6lt9����t��/p��D���q������c�����w�8�Ԭ��C	�i-���DLP7QR:e�w�TS�IK���FP�z/�'Ŋ�Ӗ�J��Rg��p��^��T��	bv܂��@���@��i�[�SM$ۿ~o˕qt���._:���=�����������=F�e0�G�	!7u�*�������/깣�gU�6qa ����=Y_���;2�AҦh#��n����#��l��j���ɟa+��q��f�gn�Ϻw|���=���ߊ�a�u֏؝�=2��lHOo�>�9눋�zֳ�o-\ﳒ���rʆ!�oa����v,�yy�e���E*�Mɟ��_5���������W^�&���P��j:���w�Bi��|%�*��
��m����-�C�w��pc&K=�bb���[�P � ����<�"��Ε���m�_�٢��gױH���g?��}���ғ:���h�KF�)����VIـ4�.W���D�.#�]��DD]��$}_`/*����|��K�Gu�0:Z&�um����ְ\�D�� >F�>p;b%@A-;;jUzũ"�����+{y�W���Q�٬Ǆ�
�2u�}c�"�b���ft�E�����+��V�'�,I6 &��A� v.�t`߃�bE"TO��lkSB�"���՗�_�h��O`����S{�z�]@Z�� �\������L��b�a��-�V�Z�[�|璓١kLE(^,����'��;�!R�!�zir�V� ��G�����6z���v���Z�8���`�ru�VvQ�?a�0,N�[+�۷u�k�J�k4�w�~�9��Ή��%��E�5��/�>9/î%ꖟ��_��%��i*ς�7!ϔ��y���y�vTa��)��3K3�«0ȭk'HUk����������. �F}Ut�E�?�{�e��1�u�$�ܣ�䘈Ѯ�>����t'��6��Z�{�PP;l��Ȩ�b�VPW��d3P���j)����p�3(��N�_�6ߎtu�xu*Z64mo���e���З���,5�b[aG�z�<���P+.�mX������6\Z����bZR���<��-̓���e�;� ��Mu���d���m&C]&�6��/�p3�Ȯ�5o��)�۞��P҉ �D����[���"C[n��Q-
��[~<�S"xL�_�e�szK�U���D֤-� ۭ'��j�&&�<>�:/�0�.N�R('��-l{�3���ٴ�o���9'�w 5����b�Mk=��p��׶��BI�vu�����x�̈́�������<�k
��M� m��!XU��u��a�|#���4����,$6CO�l���v��F��KB�Љ�7�<�r�3|S��<[oX����y������P.}X;�v!�vE7W�o[�o&��'C��ǁ��I8��-�)A<ٳ��nka;�X�`���� ����C��@�Q2�	ܟ\	)�]��� �����R��f���