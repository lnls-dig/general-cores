XlxV64EB    fa00    1ca0�?�� 2\��̢w�22��m��$։a���G�����ڑS���ұN����c�~J�U������,]����O��r�t�eh�ءW�W��{�2)cv�3� ���O�� _G�:�526�����6#W�����z��cdlj��!���k�-':
:7���Hm�AaʷT���+n�5��;r(�d�y"���t<�Ě��V]f�5®��+��(��5��ϗ0�(�@$�H1�*Q6&Q`#K��u,uHN��m��3=W�x�� !j�i�'�P��c����ׅGYÈ&qƝ�e��z�RH*�/8D
�t����_E>4t��[���G�~&�g&?\d����g'����{�S%��=m0߉�kQɪն����ޑ����Y�1�4�Q^
i�ɩ�C@�foZ.i/S6��zE&�on��Q��H#�O����lK�u�<��;��Q�4u�>e<k����߱���:��pD�����2�m�Z�dJ��#�@k��K�6��I�6+�7�ąs��E����;���u��U�Ρ�/�C#��^&���������{��s9��8tކT�S�O=����2��N6>�;O֦�Q\ua��FX�GM��3	��d7�m?Uj4r2�/��c؋=]�~B���A�6=�:�F*�|�.�"�d���2�����C�a�Gf&)����<��a����	��>,{�>�|u�k!(�mDa��Ħ��#Z,"R��TE����8 �U:y<l:	��@�!�۱v	
���&����;ff�<[	k�Q_ԏ�e���x��{�H�>����F�)���>b2���鋜lF?��H��O�׉﮼6���'�ryd������K٥�rP��m��H����k���k�Uj�P����.4 6Ɏ�O<�0^�6Pɋ�R?��"z�}���]R*G�4������[��J�u~��um�4��l_��Qb����V��[���94���N�ϝ� B8�ZC��@�V}7̲u  �4��
SД����w��d�l
�+Ę^�ز�w��>Rm��2�69iA8G�+�m��>D
Z*V�n�k��~{�?�+$!�~�ZQB=th��\܂ ?��
E	 �=Ǽ"$��F�=�^
�����޷�}u�aw��ͮIM\�)�D��%�W�~�Bk���Q�e�U�^U<K�:�jsO=�sd	�u+��'~���gec��$��3֟,҇lШ�`rPfܩ��_)Z��\޺��E��ih^u6�^y%,aak �9�Ů8'��E�BDf�f�c���d8�G��}�F�n[�\�p�!Ź�@�]s��0�dL �=��ە���lߢ���]#P��j��H�kh�_�4�x:%����/n2։�_Vu��P�����y�gbr��ؔk�xj�K,���U���-����m��S��{i\3:�9�J3�B��n:�"9G~\gl&p䖋��yYn�Y�[>����)���7 .U��p������.�gQ���hf��U&B���$2���Q�"��bɵ�q)��H�/L;[�X%<��E�:^��Z�!MJyMTh͠�W�Dx^���l���%�uk����\�`p��<�'���"�BI[m���ZK��"��hWي��SrVJW4Z�;D��ir᜶Qn��¡��[�$�����leD��xӿ���,�TDTI��Go5d�H�X�K�����L]f��Й�<�R+	ߑ���\�7xy�Õ��<x��p�ڬ2ⷁ.Jl���ԩ�j�������o�x�DM�2�ċ�̩<n\C�g#��K�a�٬l�T��hF�Q�I�¬��1��)�.D$�9�����J@F�j�EL�E{<;�)��*�����Q�J33����l����<���_�z}l4�xׄa��?U�hed�L@,[��}���I�t#By�ϒ��W������iLU����W!�":��(?c����ʱ\ �O� �Bq�Rz��V<M܏WR�O��4��ī���S.>/���,{�̿���/\�@
=W�u*y�F��A#�q���BnV�\MdQ�<��/z��	�x�A����h@�z��l�聟(s)�T�YD_�'�x��2#�,��v�;dy�'�l@��o[&�t��ū�x��~���U��1���[�\�7N	KL�X�T�`��J��URz���І��գ�c?E���õ�zIE$�wV$��a�	�u��Y�"���o	fK8w�IE��\�Ƶ�l��}+��7�B��>��v-����,��X� =C�:�:)�����2�^�9 !� �v�i���@�s��@��柎c���rz�<���2>�q�<�fzs�h�t,���:ܨ�Բ����sZ�<�_q5��l�`�Z�-��J��#���͵\���K�طj?�<��noχ��Ta"�����̃�pf�u���L)�w�<<���V��6p7ט�R04�hFLM�5�b	����Sv#{.v]��t�r2�/�:���_�H��wx�D�h�.[�d��~.vRbT̆����L���LΜ)��������@�x�ww�u��������oN�S"��m��)2�t�BŹ�Y[�n������0��/~�@(��F��;e;�#؄�����JA�X*�d�<s��`�YC����Nz�&�����$�8:�$��ֈ�S_�P�K�`!W}�PT�{G����a�5�;�2y�,������T�ޑ�o3Go�`P#P$�0X�l���i	&�w7ǒjB���FYq����\��볐|��:�Q����R���W�m22��9�g��`�ZUk1�X?l�u��>OVg�~�����c�[�w2��:���;<@W��ޱ�<d *�hP���lt4?������!#�lC�q�r��6��v��b�F��@���q
��5���T��c�/WOs����*��~x4[Q� ٠����/��@�	������D2��=�D��"8D��E�����'����	�kk�c��߉�gI�r~��c���$�~���[�:ۊ��d�r��g^�ٕ󆁹o��^G��DH�a��b����A1�2�H`z}�-��/u�(�eI0ֵ	�O�0�9`�o54��O�&h��q�����aP��F�� ](6+�Y M훥C�w�m<]u1��郃����)+o\Ĳ~��v��E�Vn�J8���R�P��� ؐ�,A�df����ⱆ��w�K鸁"ø�uK�Ӄ%�d]�f���_XBiYz�d5����w��*�Z���Yh"�]�P�ݫX&�@nH�i��� �ޅ=��#��h��M&�&��k!��;X?�: {J=u���Ɂfa�0��i����F���W�h�VL��6���+�l�b�g�R7C���Í�oJ�KA�yun�"U,*�����F����'��� �~���� 	�7z������\�����np�L��me��s��V�Qm��zH�"� R�DY�����&[e�}�@�DM	�7����ȵ
oCZ~�6Y�t!�Q����K�
3vh�o�E��I���	e�8ā
��wp�$�m��lU�qU0 ���į)
�誯��;T�
V=n�84��SIV3F�����O1Xj�s2�>�z����謶s Q�Ö���-hΉy�(r�̸[~	��PVn�4�3RV��M�R�FV��ro�.�HT��� p���Y�L\��6w>T�8�۵�-|��<��O�NZ�dGO�>�-�Yԁ@l�c���&�L{h�PɁ"�Bzl��D��	�d�#��Q������3�\b�������a��H���ݍ�䠾�q�!E������L������*�P�Z/x�����&�7�I 1|!�z
�z��ӊ��3�$Gw�n��R�n�:s7/���>��n�Z)
�`�
�r����@��i8.V��h*#��46��Ӹ���Rij{T��P5V*�ؙ�y~��<�(�A�k�'�"$B�*�[nů���k�h�9:u0c&��I*�L6�'���l�7@��0&$���8Mt�e ���᷺�E>�3�\�w(�B�S���t�6[�x�#r�����
��׺H?���u��E,�Ѐf��n�m�5(�f��o�զ��V!-���{���=��r%�����T�=Kuh��	(���Nhtw�VRc�4����,�м�����
�fR ~����Ȍm< Q�T��%4��[��Y�t����p�3�8#2��G��~-��c��@���n[��Mr8 �����R��oc�d^4�E�]
Y�t=UV�h�r�����xx*V�TkYH�D^A�k&!��=�:{�$̋����B���6z�B ck�`���n[��j�:���p\PЗ��g�N��I7"���)#�L��(�~j,QF}��^+�����hl�6�l��{��'���V��|�X���;����d������
(�ʿ�(�bտ0v��q%<��I.$������Z6��l�'�&�<כI��Ф^�F����Mk���֝���ڤ�������	_�dY�X;^����_��$nF���g�c���^���Y!�eȤM����Y�+!_����� x\���Jx��m�����cӦ���!��k�g�=�W�Pvm����u�~��Q�3Ոb�z��t�}Y� ֓����ÿQM.��� l�d#E��#v���.�$}��iv��8����8����]CE����T0���kc�;�ȉ�m���D��f�c�\���^ɸ���L��ܻ%'��ǡ7��.�*auۏ����XS�)��ۅ=@rF9{�X��o/�;a��9��%��������"T��⚠a#����H��u�څ��b�i��gìc���k��\��0:����7�>��6F�K�P�eV8��;�� �낓��%U��kdQ�vhg�,ϖ,=��C�cm���f���3����,�5��D�_�	�5���� �X�z+k��4��y·������x�Q�o�[�Y�;��i�х�K���Ie�1Z{�$�e7��x.�d���}�y�i}����/{�>��D�(E�߸g�.���"��ו��h	 {�'�?ֱչV�Q��ӑ8������RR7�VYd��i��롐�W'�nțvڭ�	��̈́|W|a��g�SE��`�>c�A���[��HA|�	K�,4����l�u�DA{�_P9C���v
˷��W�����/?H��ՎZ� �� H\�2D!�2��5~��_��(�p�����z���<��0 UЕ�[o@I]Kc��J@t���&��D���s��_�]I�� u&]̝�h�ȿ;�]��F��Uc��)�t῾�B�ᆞ���}��^eX�ܭ�s�&�9L�r�?�mM�3�nl>��r��aD�Ǖ�G�t�����c�62�U��>��P�M��~a�$19�N&:ݦ�}ry�F�4���0j�EȠ&��g��p*��j��G��cO�.�w���O��5�' o��K������@�I��2] ~�w���s���,ө���᪎ف�A��!5�I�u�"��A��'֔*�p�o.�IB��=:�t@�@n`.�c�n��qnH�eK�.�fz���g >���.��d�+S�saQ3+޶��S�?�梽�����Z�Xj�hvvj ����0�ARlL�l�!i���x<�e�-$�n*#Fa�?�m̉������s��B���I��@�I-B1�N�*�)z��j~֨X�;p)f'4���3�P0t��+m�f#��vټ>vk�k�� �7S�>���0A�0:_M�
���a8���֌�z�&��/���QV�%]�|O&��O2�{bE#�(����
F�
X��h��"�
�ɗW�^�D�obeՀ8i=7�3�7����t�i�fm��͂n9��o���v��'�g�'��Jp�}Ē�JHZev/Δp��T�V^Tx���v�ܾ�bF� =$[*-N���b�֖�膳UΖXTc��f��.P�x	 K�JpK3U(���:���Ʀ�~ ����/rL�EVU����0��+T�
��D)Dmq�|�"ҏ����/�'yj�3���\Aʮ0W8����bQ�00;�n�c��L�2Qo+V=ew��:I���˨@�Ѧ�9�:�g�oS:��6�<Қp�%[e�s/@�	$�B@�o��̈́�tVDZ:�X�u��ݚc��y���E��p1��wYmjy�"�kK�#��2?���T��	P�D>�>���An�H��]i��֎L����OejOt�;'�S��Y�S%�T;$�����4#�æ��+����I����Rk�ia�&Z^>�sL�ݚ��	$�B���	b''}���BEz8X9�k�B���Wʻ!S>=�C���U�>����B`=A���R���M_s,ߔ���uyT�H1_J:�3��&ck��L����	:k��ox������UF�a��[���7�*�O�IjH��"E�������nո0
�Q6��ȂgAL䳀����z\�&����!�N����I�3�C~k��`~PZ?d�	�)I:9@�nѭ�t1�L�π���}$��<Np�������x;H�7�\ǀu�N{^�nR��M�E値!~7�[>�y�S��χG�W��{��R� ɦ��0l���m���0Ԣ�W�s>����˥��v��F4��A��+�Z֯��F��L��ֱ�W��L�l�N֯��uCUb��*o���m�_����� �Ŵ��L������L�~��P�_h����r��f�����9	p�)������gb���X��	=�G��j	e�!�|�S��;�_}�uxZDo%�;��{�IkPgh�� ���Hy�I�Y�Q݄ֈ~�����IԶ��|��n��Þ�����o.��,�1g.{^ȤF_��#N묔�RW�������b�E��h�E%p��y<8��=��;e7��qw�{�R6�v&?C 7���1hq��	��V�˨;�I�&`eBɜ@(0Kj3��m���P�[�b������"O�:��WZT���:9F"z�E�M�C1xbBׂuD"�ֲ����+)�����W��'��s��,*U~�)YC�0�U�� N>\~�\����XlxV64EB    fa00     cf0+ΐ *�$�t�|��hy���e`�ʃ���0���b�F3��c���,���Я;�!`z1I�v
��o]*|eV�#/��oc�>d//�������C�q�|k9�	�1��q����ؾ�k}��3����`�ƥ�1�ͼ��K�����Z&�#(����/�wZ������P�'U��4~Mi��̈́��e�B��S|9[��/�.J2��%Rz(��VRZ����*_�g�<�Y@4�����f�2�R�^���a_ld�je�1E��1�)�Ť46d[x�����/��#��ձ�����V
Δ��^�	o������,�	N[�d!�$��R�QN�&�����浮�rYm����}� -�T�@�v��"Kk��BD��Y�?wM]�'�\m�f�U�#5ܠ�okcv�Pzl^����ZD��n�/iaWm�2q�ѥR�&YX`Gj���~Z�}�Q����(I��Sb|��Z�&�>|�<���Aߍ�"{Me�.|��h������¹l7�A �e���g�!�4����+ktT��;(ұ��Bq�Xd���,�eh<���-p�
>�I�*��ׯ�3O{��[d�$��L�ڦ���]�=�N���\=틓��.�6L�Q�0���̍�0�PϚ��0��Dy��	��C����Y��:��b�~��l8�����ɑ�d�{���`_��hZt>���+�捐3�1T�W��C�Mn�N���^7�v|���i#/�k��~ʀz�sך�
��)f��x�;��sG�k�\�T��d���ų@t.�a~d��WW/e˧��'h��y�ce�,�a�R�e2�O��@��vd��xx*��ᒭ���Dq�;����d
�gefnfd�=wU�C#I��r�U�S8��7�YϪ}:��'�f��.;��������	<�Ý���OT*�^WD�?�N0�R�c��U��$��F��L�;�f��g�ť�b�Ϟ��y���!�M~Ťb��v>!�>��'�b�x���xnsx�zH�UR���5��J c"���qy;��؂�C�� FT�x�7e ~�-������Z 0����D0���#�2�U0R�$x���C+��ա�>��L 2;���KN)��Z�3�,�r��D{��ͿvU��n*�{2�e����ن�>a�L�\l��[r����,���櫕[����L��g2X'.�k�Z^�ZV��O�jF0�g�ń�'�!(����9�����Gv��$b��6��j)��Ž�A��MN2��~%��Aɬ��B:$��dд��s-ł�_0v��'f��1� �^�h"0��un�,�/���2N�
���DX��(E��E1}�J�c�Pf6��f�7���+7����^���H��eԛe�&�h-g����΍cZ���7�J�&�i��&�J粪��+"\�P�������	������-�טw9��H2z��x���T��B����au]����Ų&������(�[�^��Y��M�|�r�#�n��ͥh޿^$"�2�,�d�A �qk	`��:3��1�S��Ր�L��B}b�Ur���ᮏ�[ڃP��F���ʶ=r��I=b�����&��9krO����ut��ݚ{��GsTQ�r\��� $�=��G|#�h:]��:�XZ6��ow]�qL�͎��������zDq��ǒCi;1�&k�TIUj>y��R0/�����c�SeG���e���-���om�B#��Z��&P�{�3�W�
(Hv��i�Q�Yk4��\�E���:�b��Ǭj�G���E��LT�n1����3�|��@��|���Q��݈u_q�$w~M�<DM%-���P��+Hx4'����5�i~|��H�;�������1aǡ"^��]�����r���a`t8�"�Z�PS��A�� |S��D�E$�;r��.A��#9'{X;��ˆ���T��duYs�y�{l��o���#�{
.4�·]�pi�BUD�qV���@b���ȑ�j)�����h�v4��"r��<��{}��g�p�;�߼�Y��7z��D@'V։�"3N>��8���㓎�//�nۀ�����%r��2�Y�IA��i�I�6b��
��\k�Pȶ�>`r�o]Io��lQ
�XS!�����S](h�G`c��ҿ|<Cg���x�Z2%A��Õ���U�Doi6�.��"��;��/�y� ��AS\X�s�Ϙ͓��BbXfC$/�<��܂��dH�ׇ�~TWF��h�jۨ���a���>�i��O�h+���1�2!�p,�t�XCI�:�[A��#e��'�� ������^�h�Ke_����������8})��ym�y��ґJ?���̠����fq!�����{!�7�D��,��H<�y���	'q��/�|>S��3��]�d��Y��Wy�?��h�3���PQ-B=��0���e\�9��s�=KbL�S�Gl���a�]��1*�v�sLм�V�H��������,�3i�4���I0-hY�R���v8.�����s'w.�k<��N��N����� ҦDڼ蓮ڬ��g��J�A�ZP��(7;P0GM�ۜp�>mB=Q�	���J:P��f];[�`e=������� ��M\������[{�gx���) �T�\���ޢr��y�䟣�M�#;����j�]�f�.��b'�6�1�����w�����Cǫ<e�`4>W�gw��I�%�nh�^I���׻C�u뚛D8R�E��td��  /�H����"8��
�*cc�`�+80������+gڴ��]T�P�u��V�+������q��jX�(n��;x���Ԣx�ՆZJ��ǩ(�C�n`�nM�|���qC��GhO�3L�gF���\S'Լ:�K�Z;C�,��m�H�<�a<�=Om�g� G�83�V��8����e|�"F4��qv@�#�iP�r��!�cR�ՙ��z7$P�/b���n��en��j�l����Y[�o��*��*�g�d�����:�W;�j ggZ��M����䫃�M4�4�o]"Y�f�÷��S�ƴq�Po�-U(��8p������V/?�=Qx�F�+v��D��Yb<�(�z�������NI+t9�G!�ښÐ��>�ʿΤ��\N���V�>����6<�6�ғꓹݟ����ksӰI���դJ[X���Ș���Ȑ��M� ��fr]�<��@��c���LM�F��߅@Z
)楐��XlxV64EB    3ea3     630�9��|u����(��y�y%N@���w��);ap%��GZ9�"҆5^�E��$r�+e�����^r� �2C�E%P�=U�i���/��-=��;�o�$%����a�}��:��h�J���0p\����~�7�ѐ��>ZF���[$G��}
*�MU��c�I+;ı�5V��C�Z���Awv�4q^ݲ�0F�Hz����$�G���Kӣ&����Ra'�Ah�Y{����˛#����^�z��`^��5 ��?s:]9C5!��O��oaC�EA�*�2unXy���v&(��N��MR�r�q����.��Nf�GJ8��ޭ�����-Rܜ�9� �j��͵���)ο�JոQU�G=�f�H��E;\uXY�|����:��R��|rd�D$3m<��G�!�om��� XQ=>31�|nRX70w)_ ��4���8�y�t����S��|qΔ�R�o2�8�iw�+���W8��sF��L��1#Q�{����OQf?��������Dψ`�rTw��Hӿ%�
!�2���z�P�g%�����\�g�NS{������@���>h��K��7{��4�9�fe�J�MR&G0����%����?��W�;'
bgy�׻G����ۀ�D�2�׏�m������H��_�z��,5r�a ���}�ԃ�35��z���5�Q ��,s�'ъ+�p�1�Q��5����EC��&BN�4����$�>�{c�ll�ܕ�P�����-�B�\u�bu�4S��u�dѓ4mAG�|�6��zk@�*@�~���79�ՠ�%�{-���a�7�}_�)���.�`hy�.\k�4�(�F�-�WEº�c;�FKC� F��J�Ѿ��C4��M)ڋ̇:��q|�5�f�n��O�|<t�z�@GdoD��l��˯�Jk�)�
�Y�E�x�=��sW�E�;=,��Z*��F������8�!/�%I/3�7ِ�����gw�W�v�g���Eٛt��G�̗7i�����pola���~yn�6�� �ڟc�N��U���A�d����<sKF�Ig,6�:ZA��޴R�rl5 ,���P��ǖrlFR	�Π��
\ R2���G���VC΁D=D�;4l��G�A6
zURh������7��ʿsF��2����[HnsdTC4�`���;kMg�� ���hIx��V�E�,
�+ӱ-�1�_L:]h�||�b�))Q[�S 0�r7�B�Vt�Z���25��Ӛ}<O������`��n��8X⇺���1��x�����c¦���&�
��,$��^(z֕��rE+M�	� �S�R�P-��0X���J��D/��JI�/Mi�`�]UW.h�1'�Kl!K��UsDGJ˫kB�x�TLN){π\ �{�C�,�Y:F�-gӊ|�+��vo��S	TM^�T{��[z,�
��R�N���GA�~�L7��ݨ��:� '05�0�@�V�R�Nl]��ۺ4����[���a��ZL*���W����ψAǙ�f�:�f�