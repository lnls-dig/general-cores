XlxV64EB    52f2    10a0(y���)��Bd!D�I�wqI��ݏ��2{3��g*w��O��Ll1�����{C�-����t�LnO��Vv,��-�C;���p�-t
J��m����� ��l7��k؆H�w1�������1�1 hO��,��^��e0�c��4��0m������(M�2y�����O��l�E:�`���O；��{�h=�Cb����C"3�ʕ��g)���<Z`�-kfU�u!���_7i�5Y B���z�����rWo�"LF5j��XA�L�"A�b'�4�%h_r�l�u/솪����S;�N�g�����k� )[�����VJ��V\h���m�.?8�t>wm��ۯ�3�1�Fkƴ�}f�p�q�\{�&�`����yittw���
�鰏�ϝ�]2�S��'��

��A'��P��=��5���X��7�`�_���n����G�'50}�H���6ّK_5�f�;r�TS��?�J�|K���\(XdC��{��q�Уb��Չ�x{�lת��z3*�-�
�T}��"���\SQ���贞�D�L�X3��.�L��=�����@��q�2�D5����C ڙ6[tH�x#�`m;��-�eӎ�q��'�9�/��h����t���^{{���^i���7�U��:�>��A7�z��l�[l�0;��8R�y`��X����|���Fެ��ʵE�zDlS�j����C�3�6� ��Tc��Zb*G�D�;o"sy:�Ѥ����$��-�7��\7Y�p٦�g�@@0���5D�3���7 �u�Ɋ�F��I�t�8�}�+����a�/n������i��� $�`[k=I"M��#��������|�mK&Å���q(��m�$U��\hxH&�9�'A<*�O�5B�����@��ix6�)��V���Ut�� ��;����"���-��?h��D#���rdtM#��ݡ��H��%�L��8�g���sAm�-��37q� ��HA�	���*$�o0*���	im��U�u�����i��6���7<0fuV���_�8�2+�u���Cb��G��l���QU(WCM�q%����'�2��m4p��p�P�����ԅA��=����_jk$L��X�>JX��mZ���6*��[�s*���WK ,��sY�74��:n��ɿ�����^�ؔX�8"+�~ك���|h�Zo
/ܜ��6Emh��re�ݣdi4�Z~�����ރ��q��?�Z���&�x%�s��6�!��9����]ʀs�>B�wy�Xr ��)��(0��L�s�2ה50,&䱏nu�<�-�$ F��� �1AYB[�S��.m:�-��A.��'�8��u��������o!3��6	�O4�����~9����^8 ���UJ�|�a ��]�hƵH�����T���s��A��fYf:��J�Fщ�]�?Oh`	+ �<p���|�ض^�� k�� ��Z3I2v�1S`���&�����v����Yh���$L
�y+�şX�ޘ{����|��M Y~+���l�����|&�9;Wj+2���GL�7o�E��YlB/u�B!Z�IfOK��u���ɻ�zu����36Xh����f`Z%�)z
c@F�0�>�����ƺ��T9�)�R�Z��"�o*R���m��5����$��C���3����8%я+��8P��q{�Rz�f��2�8p�U��ن�;��7%��L{q���� V���n���	UV,4�:E<@:á�xs/b̮c{�~��AT5�5���r51>&4��/w��mY]o�I5����5k'���L���I��Zn���@G;��v�7vyt��,�s.����	��B2��yI�=v����e�����J�Qȍ���1��Q�in4V���|� ��܆i��!|��o��qoM�g �F w6����"�Z7Zh�N��MP�٨��$����~�T��`l2-�&���Y���,�e�׶y�f�+2<��I��GHL�\�wj��C�}�$�a���e#�ˈg�� �g�D6�r������OZ�l��L8/h���b_�LJH����Bz�-�,�	q�jӡ.�\?�Hc��[8N:�L�A	G��1�T#d��(���V�;�E�N��@X����9Q�����M?�Θ�%E����C�B~�� lv����o��>7S!��K�=���F��[��[l�l�IM�sf�%�xt�Y��d����W���a�7E�z�Yg�'�e�@h9��>�m\n��@���$-R|�>��oVI�Ue���o'�0̆G8����a9V�p-{f�9�����[k ��f�6��S���{yj��H���i��;��*�1�!B%A��T6#����G�l�h��>�F��]%���ADݒ�]$n��%�����`5�ѿ6���TĞ�)�NH��P.�i;�)�n���ݹ?�G  �o��{�M�?V�M�ʕI����z9pȂ����v�+��Aѧ����i�� ��n�Gf�|?\G+D���&�t�5J;�1ĕÃP�L嬏�.:lb�d��I�	��("Z4�`Ϡ�S#�Km��.��H#?�0�kO���j��#�8�P|�d��1j(%���X(�����_Ո2j�6�#گa�4]W�_��q�H����83�����ǭ���'G<�0�wdכ8���k�C�R�]�K*�&2��ٓ?>ɗ��эd(�,e#�fގSŷz����JVg�la�x��WkL��[$f9�[�=��! I\������	Y[o�BBgQ�?�F��Ҭ�W-Xk����g��f%�~��_�\�I,-
%�$�L�\FtP�f�b��A�b�l�9�0��5�b2i5�=I �6h̷�'O��
�5�t�Pe����X=��+a�h{pڇ�l�?��?
sT�4c��SvA�΀���j=����c�my/}R�O���7��&�X2O&���oϟD��\�Z���;��pfud�+Ka3�X~��#�e�e���кL@��mA�H��l�H��ql���dㆅo�����!�Jgf�dv�^=I/4e��[���r�+3TT�x+��7jr���o��h�h��M�5�n���VT{�jŊ界�"��*q>G�x���F��D/�O�� ����A�Hm�u~F�yC䴎��`<����1Ҝɮ���z����:�#�*0��o��^�^:���¡X@w�ܓ��xD����6���cۡ��)��w��lpS�\*�����ƍ3�|!PO�eO�m
�yM��x��e��]s�p�1i:睦���Cz��t�=^7�T���ّ6�yoZ���i�j�_JsX2�N&�/��ݦ�hs���Ef�JG���I���O���V缠�A%�z4Er�S��#e�*F�}�<��o�`6D��]�s��?�O.`RL����N*���D��L,��{�EF�'U`�*���2��K�W����A�sRjL��!gCSuA��PN��rB�^Uz����r���G�r���۪T�p�O�����r&ؘ�[�
���ڌ�$�-��'�e��"t��E��yH��ߕ�od]��B	��(gU@���n�bbX��[�t����oñ��l7qF�$8l5����q9�\� �s0�g\��W]yį�(Ɂ�q�"b��|7Y�H��L�rk8�1���8!b3i3�s�����r��ǣ@�{WN#C�`!_܊��1�( ��>3��EX�H�1�Һ�;`[�����<�
�c࿐:�M��G���5��`��'밿M�^���?��jc�j�,W���ؚ,̹��<l(w_&�{�p{x��<c��A�����y'EB��h9��	�?D�e�~���L�#\�Yls���H�{FTWz_·3^/��%5��ǜ���d_&@�A�v3�t�����u<�2�+������_�/�l�v:[z�n��DdDc�L'���X�ǫ֩�ˡ\�W�.hg#%�B�;A��~""��ʁ�&�;e���/�id���-1�a��)xbC��<$w�p�G_����+�!p1��t�	j�'�_nq���,~�)������=��q2:���v��#t��]S��(���y]:��z'���u�c���kL*e:�݋�͔�X8��Rk�z�Ɠ�F����W���E$nBП���l'r't�@;�����U�Dj�jO2�