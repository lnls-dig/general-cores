XlxV64EB    6ef1    19d0�N��5�7�U'C�Gjr	ppJ�}��!��"�\w�h�,F�N��GW�|�ϓf��]�-�붩^��	Xt���V����o^O�=��ϵ�"3q�e.�9�F�	-2���%�68��ꏚPA�鈩?fh���zM��]�f���Mk.U�E2�GU�Y�덴��<ȿ�|kL�ѩ��=��$Jo5�L�;fڈ�=���*0�̕�pdZ�
�Y�����BH��_�Qu�w*1	z�:e������4�&-=T�֡���V�{���7?X8���k�%�7�Fڤک,��cO`/�<-ᥰ@Go�|,�6�o5��$a�	z��8�6Pn�%�$����'��-��k"�+R�R�<�]ȩ�<D�/�0
�>V�d�hU��"b��H��U��Sf*y��AP�S��#�*K�w��ߕ@���-�������X�'X�K�1��<2�tg�_�U)�鱫���H�︹�׈���XĆaR�%��D�a!���ú�J��W\�7�y�6ݛ�\�bZ��:;:f~e���j�0c��a ����җz��:�7	��EO��9�L|���P
� ��P��G���r,sݰ))����l��D��$����G،�]�~K��-��z1��=T��si�&��X 2R�R�h:l�����v���������}.�xi5�#d���]�\��k���v�x��*1F@��������"f�{�L��ߔK�c;+u&�Q&#�l� w��7ko�M:�/�s5i��֥��?@�y�X���LޓUv�$���q}� K����>\���P�������|+�W�Hn�l�c����|�m�U�%^�eV��dˍe4�?/4�ؿ?+M��-]�z����S�ef鑼
���%����y��H�C�OǛ����a鋱�JVc4��~R@R�����4�Got)㗐���Ͷ�d�MTd�9��H�NWޠ���~j�jj�4t 	CL��; ��b�&t٬u�[nt� �
΃LAS� �h�.��Uxַz�
 ��P��7>�����}f��`p������<~Z�z�(���ݣ��/�؊E�:3I%�
��?
��ߙ%��\��]&�/�/+�D���,h��'�����/����!$a>��2L�)���D�o��R���PJ��}�@}�W1h�c_=�Dr�M~�<TkɋyX��VW*�IR���oP�	�G� �1|Q֥191�7m4�&����:����>2����D�M*�2��R?d���X���=��0��:o��i�%��x�������'{�:�?���ά�� zҢ��i��/�=����a,�S���܅{"^�_va M�Y艱Q��i�:�,�a��E򼫇��i�-8�<(���ߛ�,-<���q��zV�	�D4�8�B�����v8Z2ɮ��TѱK��aU� G��"ɒ(	.�N[!�T%�;'ۍ�����][�eW�ߝ�i�4�̷$G88�
��M�	��9}�S�(������h��b�=�U�@0��	�*�uD���Ԫ�_#����ȶ��'����=	|��+�0	Ub��#�{��Rqk�!-(���i#D���E�u�'�	��L����k��w��R�&�b�%�%��͚�q��E�V)�V�Vp����h7'.OL�����<�^ &�����[��^1�Q����۝9鏪�����E�g��=
Ş.v����z�RK�ڬ3���5���O���S�`���<��xtBܽq�%����CT���錺#xy�=W��b�aR?e�b� �z	�EB� @*MR�>f0ڠ����>j�4��׷,񮂗#�ؼk����X{�^�i�(��W��`��Σ����w})g;����M����H���L��
X�����;�i�ߚ5��!��*O?���E+a0"o0	d���M�M�[{��+)@([����7�Y3r�2����SPc+;=l
^6�0�ʫ�	&F7 kE?ÿ/���������p9񖈓�ޖL+)-�3Bm���S���)S�\Y)NӺo�{��"KV{sE��!(��x5��g��~��0���p��D<Q�<��LG8�-�V1�
��3H�:I w�D=��ܽ@��Y"����*Ν>����D���N��<�2��Ðh[�>�Ĭ]�с>��?:�{`�u/��x{㸷Mi4�_?�p�QZ�	Q $bl6u��.9�4� ��E��a.��Pܫ�wlW����6:%߇U�3��!�#����`��&�7�O�d���(٥�Z���$����+I#|00�� �pB�[����k����@��⯧�;��+��~j+q�R���\�����XQ6�=��4Nx��`�N��~��m�3�C�]���	�5W'�+u��)E��Rc�e��QBR�z�SQk�g�Q��_�k�{w����v��1"ԮT ��*/��2.G��8w���|u� ��D���<a�.����k�Jb��њ�9�9��)���z�拐]�����F�֩��ʹ�B�aH��,��b�[�[ҫ
#/�Z�����61I������YR�������
Y�������}n���ާ�"���&��;��@`����$L1�jH%zR;�QZ;�o�e?�|�W)�|P$�=Y]h�M7��}8C�'�]5a�c����z�3�H�~λ����e߀k`G����w9����v����D�w,�~3�^����ۜ�s�p�@4o��]Nc�"�"���ŕ6�a��/�nmv�o:�50�F�h�2�@��bN����e�D�T�{�>u�d�#��2�R���ϰ�=T�0� ���l���Y�9�۲w��¾��.AJ-�R��o֨�@2����xJ�A�;;2Bt�6�fA"�-Æ��[ �d�A�ouW�7�;�y�цCrY�o�R��eV��#���S�8L9CG��0^�+/�(����v�����A֪3N��y�d��X����Eak�H���0�=��B���Ʋ�J؜�Aa�`K5#��~	��@N�!�09�`<����S.B*�� (*�^#ѲY��q}� �P��� �� P�N\)@
�p�0oW������*�Q�� .	���j":�q�֖��5%�vM���>Mm��818�E�S�e$9@�LOYвj����>��p��������9�Б���P���8p�3P�ޗ�ߛh�b���.B��8��e
�OO���K��@w��i��
���A�$*2#/�c�qɁ��%'�<�Q���W�?�2�r�����9�BX���*��e;�	�_���k���5�܊�ڧ1T٬
��m�
�_����O���l����M� ��$�)Zс�P̌���b>�Z����=QsR[E+����ʱ�����\�(3g=�f�m#�ѯ�|�������e�&�8R���V��F�/��7���QQ�e�?Vk��k��xΡ�O�䃠���0��M�l������V";�	֌�!���p�G`,�Z������'	݋�	&�z7F����#/`�qp��h�A�n��x}dM����ԑ���_��`�`�'���96��O�ʚD��SA�D�'(�|�ݏM<]	�J1��=�6A�.Z����	p����5_[�uG�#�����yV��Q+�4Nk>�1,v�@��[�{I���l�}-C�d��c	vD����3�����y //:X�;r|���;&�UZub듇I*[�B�_/j�6�P+th��} �u�S�F��t���@\/@$[�C�m�3�����{���|/�l2��y��fixZU�n�b�_~�������~��/�Z���a�>;m�N�� ��^#rKʏ.-�(j'e�����*5�t�B�C1��h���4�ZWU��0���
��l<XFT�稴׳M_nzmb��M���3"�������[�]R���C5�Aa~��z~7��w� �q�M�A�P�D?����|ty�w���f��ǫ��52�#�Z��]�p��n���\U(�����%v�ZmLS��>��ZW�%��M�Da B_��B��V���������?��n�!�'1����	�q��� ��z�Xn���1��aK��}ܖjg���V1�v����G�97��+�Џ�����M��^�Z�N��9��X����h��,�Θ��3ggl<�K��<m{BA��t�O<��D-�Q�N��خo�ch��Ł�nYx��c��wf��y����ef����㥉>M��/�����tLzˑ��8�5��?��p�
����I�s�<y4�h�ob��/N���Wd��*u;u������p��=�0�����1/(Z�v�߯$ozm������6���TџV�L�?�ᴘ�����+�\�������ҡ����z�Ľ�Oˉ���>�uҩ/��U���8��A�X�I׶�/|\�-��~F��p���/V����ӆ���[X��Ҫ��T�^�p����S6%���۝�Ͳ�4m+�r[�9D��1��Ia�*�����ڒ����ti9�P�/��+q9,��J�J�ݏ��8�!�b��X�{�pLs�n:�Ԇ?N��|�� ���Z!�]D$�k�yp�$jF4��̉F�R�j���f��^�^����œ?��=/����:��� v|�^���#:,�.6I�{�^��ΒR�DJ?�y8S!�e�������֑�
�|��C]Ɋ�{�kxk�Cfm~e��a3kI���Gf�?T��Z��Z�'��]�	���A�8��?&����n��6�w�O͏�I��╅��+��R�~0¨�dl���Z��gP�Q���z��44�T:D�(:R��ϨO,�qԝ�w٦w(��\�l��X=����h�t�@�I�|$4޲d�d�PL�\�q�C�/Q��6�yU��s5q٣���3���ic'ZG:؟`���PF��j�" 'l�;�H�s
�d�ȥK��V�����u�~JDZ[;
�ڲ�&~Hߺ��-�}���bIN��4_����"�s���tB����[ӓ�,���N��f�h�ʛ�E��t��z]�����b�0������k��݆Ø�I�6uVL�"���.�����!,8HRo��1�_��<7�^�,
�jb�6S���y�f&!fNr���0^�z�����Iv�&�{�i�
��a'�q{�(3��+Eb�m��&��?��sM��7���be���>�eʷ����pk��i$ ﬓy{U!���[��d�ƅ�Y2}��*�J֍�v�a��_3����!��1�<$r*��IݞN�Ӓ���)	�lU�����&��4kTC)V��8���4E��8��YP[O�pT�;�J��#2�IX����+H�B\wlF�H�$<�8����B�:�n0;=!>LO��ݽI��c����R��6�G�m'3H�Q�t�|��@��m�p��U��G��F�����A`x�_��.�ũ��/B��.X��lո+�<�zL�Ĵ:��%�.��4*��B6�_����֝��=TK�$j�飽H���F�	��p���?
@�9x� 0�7�t�B���p��(&�#2�L����xNI -�\���[�3�j`̯�7�@�=�c031�ć�(�I�;��C�F��h��x�q�o��@\L(��������cZr7�W�tG>2t��Oͥ��0�ʝ��x)�AC��^j|]��	t�v%G���'�����c����˨q�/�ߧxj#���ZG�_����g
t���6j�Q^�������L�w�:C/A�������D[��W���/ �7h��Lo�4��[��Y�^N�A53� ��]�9ßR�Jw-�D�7)�7��5@V)3�����|�k�ڻJx��P�$���m	T (J�;���Ǖ�	3�\�5�ё8����:���D�8IO�F��V��颂�>�"D�{��;�:��?�'�'�G��]�_���G�H���!\��$�2�X@�hB�o\�"�ʇoԚ���/
Љ��!���t"��@���v�4d�U뛠t��_	����E{q
� ���~k���΢�w#E��x
�%bTH�P��r������]#��� �֜6����Q\!��X�r&��x�i�4�C$�D	OzK2�D3*<ꎮ��
�<i��#��K��T)�y_h|�#4 V���\>�"i`�Y����|�*Sy9*Q��*��@ؾ�{s��)�k�J�V-�TF�;[5-���dA�
��r׺�U��1H�u��bL���G3��7i��֓�s�����~ڀ_<w�~�NH����� �.���6�8p�alS��V���!P_�HJO��u`h�B�E���,�i)������/
���[? ������@��B`"�)��S�$��&'Я'�w�, j&�����]a��5�