XlxV64EB    3fd3     f909����t�nbPC�J\�-����О黽S_��_x��4�+�L��������^`�h � �:��(��L����z���pdQ�݇�a���e\��չ�W��?E��j�}^A�oo4F\0�������s���7<(W�k������w�&+�I�)xS^m�k���!��^$̨���?4�
�]�M�L��Wؑ�$$���Cp:L!E^�NX}\�����=�H���X8:~��+/ "d�rֺ����GS�:=dXe%m/3�)�j%d�v&_x���M�0!<BK��2L�f��^�2�!k�����<�B�#,�B�9o����C`c�	�LD��`g2��4�
�u�$���#	s���YT_�j?$Zuoi�!O������i�6M2�>�}Ni.��I��@���<�+�sy��7��_W#�ꚮ�]8f��3�hX�|��05A�4`�&��';��k��[|��.�0����#}��P����$� ~Ϋirt"ύ��iǨ����I]�KN���/�"T�^�¿hٯnҸ���)g��[n��g�7�q�+^6�8qv$Ъ͑�)�NAkg�㽑��e
Ğ�_��=�?d5g��Z6z����v|TJ�~�s� �cO�J{���ӽh����U��I|h�RZX^�`�d	o	���ZXl�����mOQ�*�}��n�Oh�&�ȅ�1s�Q�cS\m��k��@��Ȗ��-��ȋ�VX���
�����h� ��:A5DJ
���2��u࣮����⪨�]�B�r#�i���71ҕ�oobރ ����.{���B��*4k�QvP���R�{RkL�P���
�>�&':���#�r	�F͸�ˊ�g��5}K ����$���оrI|��N�u�X� ��7R|K}�?��P�t��τ�U���<�^[�<�?��w���݁(xLyDD��K ��-�:���T�K��A)�w���O_�����hs�03 _�C�������+ ��wH�B2�*��AR��Jk���S��!˸�����(��b#�&�}�e��xZ�m��!��8����K!�z!Y��:��%Ɠ��Vd��m�&9����M�+�A㸜n��ؔi��2R�9f��'�8[�݇�[�ɺF?�܋.tp�.ԍ]�Y��W�����Sa2(}W�DC������s��2>g��q�.!O��(x�����UE�.�����l�6As+���
6!X�@��`�[_�~���}��ygV  ��r��ƶ�����%���髋��&���hB��ǶF��x�D�@�bp��fݻprr�g�⹰����ȅ�dM����t �,�c ��s	�^����/��rހ�	��q;���$�Q鱚A�{�!o=!�������w�H`�Ñ+��{������{E��T�=吤����[р^fek�0���Y��((�ͽ��)f�M�K�3�G.�Vt�T�.��`q����ܭ�i��M���%��u�;#S�ڗ ��V�����z��1�?Ⱥ�=���Q�Q
��k��Ͼ���g��&g�4_4m��сwK�fV��&&��(��4Š�ep���7Ws�MAi�)H��S�T�NxO����g�pt�5f�-��n�[�S5�n;����`DH�
4��A�%����������i�D�z�:0=�|�lM^.qy���c�qnW��m ;F�ٜ�����#���&V�Ϋ#?r)ź����_5MФ"}R�"�v�u�j
@4Vid�wư��^������2��^�iL@�p��sC.�B`�MbX�d�6�kfF�YC��H��Ƿ�YH ��PIH��� ﴕ\��X����},l�n�%\�ǲ�����d��_Ar�E��t���7P�$X�ؗ �ʮm"�2��Ҵ6@BA�6Z�Y�����<��R�1��쳾�.��0,��N��^�p��25�;�$�رjq۹{_�����;|�;c�i���~!z-*�z`殚���ʣV~��H��pS��d�ʎ��$�8zg�颧�%��&�~������`' 
�!��va�a*�ãI�<kj[k��.�1pM��*�I��dS@���Q�g��A�zC���E^~#��SB��p/�p�A��{��^���!F�@ֲ��)�DW�p�o�����~�ՙ8M����R�J��Ͼ��uI�$X��·W�q2��w(|���G�k ����N�D��iʆr��oz����+���iX�K;b���|dP��!+;���BR�0�<'��|�t��u�QI���8��>tid�ߜbo���;�(|�S����;_^���/��^��[�����a����dq%9=�Y��w�!/D��ԫ|�2RKY�5�ih�ϋn�s m_�����o)�DQ|�lS¦��Й����@�\�$��F˲^Q�3)���c��*�7\C��{o��,(���Rq�A�0Y���G3�X(��q��6�6կw�� #��0>���Ke����Au��wv�ϴƿ��v OP[��$�"i��uL���i�t�K���duـ�4�6�Z��}Z 6k��c�.�T��>�A�D=��d^�$M�hS���GV�`���s�N�Wm�A\X��9���3��k'd��al|CwZ�"�-�*���� 8����0m�%MNQls���h�0!G\��ț=�giJ��
U���^���A��Wg���L9C9�^�.�Z8�ѯ{x�nDx���*���\9� m����?�̑�bc�-A�������֢V�*���V�*�/�`�f�����M�1
0�	�}U�(�}1�ƫO���JL�<������"<d<^$�?�'�Q$֝���G�׿�;c���I
��%����	�%��"7�o ���C�����_n�c��	�<�ڿ�dB�Yt2՞�6��\�1�ve~���r�$S����,Z�qɕu����������0"7�o��:c��A�����ihL=�>Cwp����{������6j���.��н�)U��$��T���Z�!mP '7k�%RL�Ӟ��Vp?� Ң��}���Fg�����B�x���c:3ֈY�C������F�f']%�Y���Y�6EX���PX5w�q�AU��G���ލ�/��_,���*��`*l7����(�)����7�?֩���`m�:�E��u��fwMr����+��E�pY_�B���X��D�l��͍���{fG=r�kL< ���,>�Z�ƌ
�o�A�p�g1h�9�9��.h�N)�5�,���#jA��P�X��s�p�/
�܈#-z�P�J1�vϯ<��s�)��rP�-?#�j�8ixC��m���/t�1���@S�i\�[=�3��+�4��Ox����1�m�KPꉙ׵g6S�*��X)��=�/g�l-��4l+DB���װ�"��I^�����5$]z�V��ҋ#�/�<����b��j7
[W|X��C�ԛ�BG��ǰ�����\��Y� ��"�3É侻�������9Ah860)�f��v+�œ���x.�o��r�f&ky������"�x��������N��?��ֻI�Y)��k��Q�j�f��}����ڂh�4��qZ'�0�@���&�H�K~	E��2�����?���h��c 4P��0�Nx:��Zw�\7�㥄$�jnsϷL�5bWq�B�0
��j޿�@g�Ns������o;��|��Bw+i�7a"�{Q>�]��EH���\�����v��&�G[-6cZ�S��~����#�_\!qF�G>L�������0*�>���/T0L$�=E��e�r���I`��~R�+M"m���u���d�����y��-#:'��d�{����	�`��C