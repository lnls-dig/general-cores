XlxV64EB    1ccc     910��?�^��I!]ݐS�e)qWk��Ȳ��ni�F��/~pY {���"Է��w;��	H*t�ذD�e>)��uim0����8 `3��O�4RT���]���'"��#���$� R`�p?�����a����,̟��I��\����0a`I��.�֟E�+�ާz�����(#]�_rټ<2kڸorZLCo	�%4*Z|��?!A�/�k
}����Ag|��+��>f�yǱ4-z Lt�+eF4N�Z���t�Z���k�4�B����I�eM��J����zs�����|���S�w�-�q}�8+-��Qe���r�c��D]Ÿ��ĭ�n���$����'������Ŧ}ԅ���Sv���<ф���<j�P�#ұ��V�m�9~ ��P�3S���Wz� iţ=)�y|��t�]�J?Yб�����*��l�!c���T�TP^�2 _�Q���-��ebWs]�H�Y��V�����w�5OP��0��v�Aٓ�BpH�ձnO�)��dD��x��鎱\������F~\�u�]�;ú�͢�=Us��_z�y��ok)"�W�oV�l�3.5��H��Re�H:��U������_3����aLo�aB�+Cz�}��i�j=ӧYJ;e���ws��Q�OL��w��|I�:4���GK򣏁'N���q���i�A�{�my��kh��c��Nr�hU������;��늚�f��i	h�m�3A��*��J�(�*�=�`r:���吹s���O�t�t�)�yq�!�Z`g��j���b-₥JfX�X�������a��mK�BٚoV��ć�T�k��h�x�C̙��b��(�0�r�����*�bJ7�k�9wJ�a�b��ykLs��  Ɔ�+��n{�L4��=(��wy���A?�ʽ��-N=8�#}о�G�k�F�\>}�V{�S�j��,D����炌R��ᾄs�a$ef��bا�{�*�����\䤋\�C@Y�MjO�>�!^���1ss����t����e{�S�"@8 N��F����G��K'�P������~r���m9�һf3���^�b9�O�L�:�)�J�Uyr�TY|23�`	r�K����Qj�E*ǣvA�%+��������&
�|A�2��e���� N��v�[�w�+�����F�<>��Z�SD����At���V^�@�}.5�t1�*T;|Ԋ�+��dK

��ggۿ�	���������i�`�p�������me�u�|�YW���"�U�ƳAS)�&W�����4	;z)w�F�M�v�q,���bk�z%M���'�z�&�q�B�򿘖�]k���'�&�B�K!*'1�?��d����_YdP����~�N�A����tLG�K��D�*�����ذ����6q.6��!�Pٵ�3m�V�)nYF�H��e�@�jq^�-?R���z�o�����o7�,',���[�F:�)l	t�K��x;x��Ri�u�d��
̈́->_��j_q�#���f6��2٠�b̔#6��!L͓���v�,���/���W�����a�rI9��_�FO��:�$,77%�E/�t/Tq�wG��������o����/	Y�\�"~F:N��1T���/��T6�
<A����l�)���_^�b̝ h"����IFj��C��&Eq��s7 �A�����r��$?�5�\.g�#�i�h%��R�o��6��҇��-��`�+�޶�ƭ�,
��>�
�%���i�����&w�X ��Q0J��R��y	Ba���õ����i�D��~��A�6/�WE�˨��,da������k���2\y�յ�-��N
��<�����R�ѱaSl�t���ӏ/.�
���QN��?��!���J�쿹z�;L=�]#��b�yD2��[�{�%�@9u��v�'��
V3OqR�sډ�$MX�Z=�i-*E���E�ĝm' �xy��6~Nͥ�]8C@F�z�0$V�[�jϥ�w�^bRN��Fg!P���*K

��F���13{�ܭ 7hh5����>n��y=\8�^�ծ�z��H��󆢱Y~>��DB�.��o�$���7hE����ܽ�� ��ǽY8�R~4�4cO����v�����F�x~�x��!�ը���(��k�_׊�b��q���h,EZ3�2T;;ONJt%ڞ��k��V-��Q��TLi�Cf_��O�l���������F�>�w�