XlxV64EB    dfa5    2a90��&S�u�l��}��,�;�S��4{���'���U��F늽I��ng���Q�W�Vp�H��Bݒ�)�`�+&4�� j��qJ-�ׄ�Z��%��5�����
^�y�dGn��b�RS�'#H�83�E��Q��b6-�`Q��3� �" [G�< A��9ߡ�v�����V�.��CH9��.{�Uq�]E�*�=�A��O��<Nϣ���3�ǜ`Kv�N�W>��>˭���p�{��Z� ���M��x/�ƻvl�@A�;ֱp�0�vv(��M>?PD,t���>|�.@�h�I�o�S-��Mq+���p=i�jE|�p��$N`�8��C烙���l��c�����7r0 �Ӆ��RP�)6(��� ;?�I��H��f�YS�("��lr���Rl�2��W�SZ���ԥ,�^3�ӈ����@m'����>V��qvW�aV���q�=/uX-?։'f6�I,��Z/�Z��+X[ �9���L��4��NSΩ ��sn ����|��pO�0��)9E��~t{70�\qC���*�LSn����wR�.�p��� �.13޻����J�ߠ�+w�3�_ �$��=�J�5O�I�6~�2�/�l����;����4@v��╀��[<��6���D/Ò���<���v�%)LA���W�8�A����\��HΏ3��s7�&����_�G�'�\�6��Ø��N�,\T"��._$% #w�4N����V�1Ɗ*���/�`)�_��\���߬�)3��ݘ�%Nl��� -1����,9Ws�ޟ��E����*��3}�-lI<5P[��>�S�vڑ9����f+Z�	��	�'l`P����.��Gs���������8��S
r�k7z��\�r '�޴P@���F���F�O����l}�+;�-��g��*���ԯc���D����G���xk�)cZ�ǂ��`@���q�՛q��)
����>���S���*��H
�z�'���S����� �k�N2^~4I��tj���k[�������w�h�}b>�$���G����t���e�����jf�.�z�fxw�𬵭k�>4�9��.�{��I��'��Wk�bef���c�/N��X悡q=Lh�#)a@�}��{���e=�{vC*���T�9d�R�5"�(��y�l"�6�e��B��������,�M�0�Cs��I�cr�p,dM)�[�"���ﱅ0r �:����-��n�e���p�n0CP�N���$�(wN�eA���ז���g �t��+���3z`�ǲ��}�>����Zudh��Ae��pֵ�z6u0���d�M���^w��6���������v� 9E�߳�lb�l���T�\�X�`�M��9�{	M��"�\SX�72�K>�͞���zĹ�L��xEXQ5����u!�[q4��z��x/a���Ӭ"�aC����
���S��
�7��+�4h��!��^���BvЬ�T�����܈0�ֺZ����4�A���5�>�QP���ɃY��:7��n4�Q�9Pn$&k�'�}LI��v:���x�i��z �_���H���厶g����m�* ߌ��ש�u���+��ԇ�Ӽ((1����c��&6��	���]�Ӗ��3�oߐ*�B�U ���O ��Z��3�ꦯȲcj�-Y�#�Cn�=M=C(�I���W��K�^�-�fs�n�(ܯ��(BI"�����vL.1_i`��l�isW�~�Z@���ּ\d3������ D*a�4�:���ƛ��F��BO�}%��ha����X�(��-ޒ��U��Ԑ 1#'J:��N�zJ�y�	�<C��!��Go4~}���s$�����C�#�T��K����6|�< lg ٨6���Q||h�[ZZ�7�>?�
M,�b 5$E�]��r  �V�O�X����#��ؔ�Xy�7�FFt.CF;��偾7c���
!����rd�m����#ELP�e��YIq�p� �����~��g�X��u|���x ��D�(��+�����i��-B���ۉQ�Z�At���+F��4�v�����~˰\�Cڡ�ZiP�a�|T�_0,V�<���p�
o��Ȃ��:��t����w��Wq*e}�Zⷞa�� 䴖�5���������+�*�.	�5%;*�����7�&��,�6m !H�Ȼ�f�����=;v��͠��i��Xp�(�tu!
f�!K�a���j����|�Rʑyή�hs�#C���ꜨQ�����g��*Q��+=�g�����:!x-#���*�mR�:^,�>����qγ�qP���V?)u�/�\�C�3��~W{?��d6��l䴱7�9bӚ�I}K�[�����o:�f��n�P11cU������Y����.@�E�S���[�,*��pW�M���<:�̝Hd,��X~G��B|�Zܽ@�+��u{�5���.�Z�.�&[!��>n�5L���9��X�)��R;j�0�W;S��Ko�`fjED�Sk+S��~�W�=���<.h�l��ʭz��M{)|�A��;��x�vu̓X�N��afK~x�8�q<D!��Y\6()�M�Vms3|YQ#2���Z��؄K��̗�v�L�umv��.�K��l݆B��(�2H�����<#��Dp^�I��)z�i����&M�0�OO��1��>���2������l�!��
��k��!�^7���3�c��-+N���B�4t#����Y��;�ܯ���}*��Q�Vlגּ@��ټ�'u�.�62٦]ï���-��Ss�\�~\Zޗֹ����9�ݍ�W<Y*E,�s���9��R��j
o��a��W�ɴ3�u`��C�0[�]�E�����&��7-��CpV}F1����*XՕ��ؐ:�������6�{���t�V�qB��Z/���goet����<�Q��"V�����L�E+<���K���n��������$ڷ���F�SS-������p��,�!��1����#k��h�_�ԒM@!G�aL"��jv�]2�7ᴢ�����R�2��`݌mQ�z9x�������ލ���(�B{�&�Q�QF��d -��/ ���?+�,����̧�b,��U2)�������-���ZG�f.��V���`�4���"�3(�	�Dg��i=�ϛ���Z6?!�]�DH�vA��XXغvb6��wɂF�aظ�c0pߟЃ.�Uk]������%��J�4����Ǫm#*;+�KS�/�E�I����� ���g�~	}�T�i���k���r��������⋑�] �J�k�����4]�?#��Wg����Ayߒ�E1륫���2�%�~�%��v <ԕp��	?�j�2k�n@w?���Mg�(�ųz����]��5������a������ԾփM�U��8~�v�9�̛��tQ��{t�3Ť'ӷ���Ƨ�!ɷ�8���bR0���U���4�䷊��uk},U�$�.#n]�D���w"q��:�V���?�?�����m=�I�!��އѸʨ��C0���ݘv�H�b�1+f�	�Ƹaj+���k�>Bfq7��� H9{�.����Y��Y.t��2�{v ���/�3�bK�C�	�.u��r`�����,��p2��\��c��u�2���B-�X��{����3��f�Y��bi�*�Y^�����D�ԒD5؁��e=�X���U6E��$,8�iꚱUʲ>�A���W�ٲ<�M���B<�HrKm-x�S8E���)�35���`�̚z\����A���
�r ,9#�&��a�i*~�By	)���B�@o<�#��o݇���`Z��*Cu����dv*+7��,��� �֖ͭ1���ND������Ѳw�A8gxك�W�5Ub ��=���6�|Wú7��I|��X��c�S������9 �eW{r�kp|��I(�����u���T  E�Z�W�&��_��f	�����^���9�Tt�v7�\���	�L;Z��qXa�\�[�yU�ʹ�d�2��	HZ\�V}�U����.Ċp�ˡ���d{�V����P,� �C���F��ݭ���T�]��@�m��Z�oq���r��~�Snuu���x��!n���"��e�Nإ�(�ii�S-F�.��pW���Җ9b4?V�Sc�֯5m�PY����X�R3�mmd�j�*nb��p�T��_a�J����l�n=��JA�ojT�w��UpY�(��2��[I�G���m"BX[)a�-o6G��"DJ����U�v)�r��7����X��v��y{%7���i|_Y���5A+�U(��b˯�����,]�<'��{x�39@Y�����,~�l�K6�JMZ)��Dhgb	@�;�D0���:�����}��F�����n�OO��E��+}$aO�N tH��R���4���i�s@���V
�nj����`�b�7������+�v�z�ҿ�PTt훎��I��S��}��[�A�ʑ �7r��l��9��9)�Ps>_�'@N�K)$�����R)�R��u���Jt��dt�z�0�0�<�*=Z��O�Η���R��#���R������f/Ļ���N��� ��1R�ݳ��#����#�r��WV��Vɨ�g����WH��C$�r|N���������z���[��K�3����t��p��*l'"��1�'6Ĳt0o�>���:�����b٧��%��f;lr���HY�O��'s,����:ف�KvHr[O�iw!��Sh�ѝ��M��s� �N�8��M��GNҧn��]�J�{Ē:��n�8i@�ܯ�P��4����E���yr�\�����\��=A��4M��*� ����ߑjsA�)5r�{�>�H�������Bu�q�8�W�a8e��\�i}Mux�����'��I�V��|� \,�}A,N��"�1���ߕ[6+�e�`�іU)'e�~�ۍee԰N�<�9�g���7.��R�;cR`�O��OCQ��N�$T�β���˖�j5ZeJǹ3�� ���ם����i2�K�S���ݛ�U�j���R��r�ST6O��_3�-�@�*���'�n��ف�Oh#�Wx3��F^W�_P@>N̺|��R[Z�k���'�Hё`���"�����myT�髧gK:�Խ0��:,�7�]�>u�{�$vn`��$��D�&K�Kghɛ�%�{�W���#]�����#i"�5��2 ��0��}'I���Ʊ0�&����o-�5��X��_�f ��`9���7�Lf�97��B;�7Uc���+��0G�m�%�\⩹'�&��;��L��){�ϩS�8� �'�w�;w�F�3���w������.0�݇pX49����ZQ
pwaw�LP��i��`3�h��J9BU�l[��(��.B�7���8�~���U���
8uj�d��>�P��f݀��ħ�3|��Y��/I�^�-9'҂�m˱��B#��+Bާ*�2�|T3����o.����l��S�?�)��v�	� ,�� �yH�S�LuD��o�	C59D���,EWu�[�䰇��;�Z+@g�58M�4픏�Ưr�%�_�i *.'� �o �7��ص���Xc���nS��G٬�Ys_@������^z�i5�!qOW3��8\�}-ˡ/�ϩxy-6�)������X2T��$��A�\pߠ�Ffќ)� �x�̔������!P^8np����c2����]C�X���l�
?N>F����-@Y� ����lU�Oe=�(+�j�4�3I���j�owcc�݌k��
�	��٘V���o������I��q�ԉj���B8��L-)䏈�f
êf��85�]�?�dɎS���}�ZF]���b�c��fgW�_�8��?� ��'=ͬ��b�F�q��g�n���Z��Xʏ� �D��0���W������v7x5�'��$pN�HB�q��t<\��=����r���
M`�T u�WE&���PY8�"�Τ��X^��g�2�Γ����P��$<���� �D�O��j�Q1R
D������orxPL��J'@G������}����\*T�c�o~�T�ԢH+ʐ��p�fA�\�T�����,���`螱Ɇ����e_3R�ߏ��*�w�s��~@��4�l,S3J�
`Q�<_�JOOH��Xq�N��&�݆;>��Tk�E���w�c6H��ގ�Df�^�bMR���<&n�Q+�Mj�mU�0�? �i��iZF��1������ځè�p���d�o��Ú0�,�A,���q�74����p��I69%AX�!��p��^.n(�hI�33��͡�WF���o���+[\��%nEȺ
7ZE���e����B�Vi���{cV,e�� �]���S���~����~��mAQ�3�����@�:�^���.��[�~��M������\����w:L����<`7�����8)>�{W��4��Fũ�_�N�ˡ�_ ���нgtBL�+>�
��=�������xɤ���N���m�,��c0��@�I�C�x�
�m���t ���`�އ9��VQ%��X6��WŅSK����'�_�~�K%`T2�v@�$E�m,u�fI����O�����iv3�Ƙ��V�^�Y��{ 
�{��p��#82����.��@�_�wR�R�=:8�_�+J}|ڄu����M������"�X�@�V��L��'��Q��kHs5%I�6δ��Gݽ߼�b�.�*�� @�k���@�KK�'n������q��9��G�S�@
X��ho���c���e��n%|XՕZ�����x�v��m5i	�>&+bq#�Ao?�&na�Ѱ�74�����5�Z`<���l617�x�#/#-	P�f�H��h!.ԨȚK,�ʻ�(�"�r��h��bV�/{�|x����J����H�^�_?E����s�(U� t���X��P'��7���4l��_%��́�>\ժ���L��DY�Z���TqN��O�6�uGI�n�/��7��p�.� �������Z=�g����\wg�#���?h�D/_�J=gs<�Ⱦp2�s�ޗ-J�A��y1��m�%��9,��}����#M�u��o��pudŏx���:\�X���n�pW���?e�KpmJG�u���?��f��;��6)� c]du�;b`tuZB���`�'��"ͩ���㑥;
�=]�y{p�"C�٪�?ncftI�c9@ooMH�%�������6%`�{��cg�t�p&͖��bL)�KQ'�7�r#���j��M8�-K��m��o���]\(��k��CN�%��g꒟eyMJl �"ŷ��&#z��+_�(���p�����Es�<B�>;����$>,j�/��~cQ�s�K�r;�c{C¥�=}HP�O�Rk��R��6�~"	,�Y(&�>}L���hɝ��V;߁�#i�,��8�AD�|��`��i��x�O�n�ERh��C�Q��9���^$��1��me���eI?�o�����J!SZ�a!�D�����W@X�Z3����1Cf�� g�Dɪ������r��JN�8����C�#�LdsS#���,����d���j�RZ�ѨA�If6�U{P�TthΡj���:����^��	!-��)��?�w�;��7�%�+7�Yu��"���)�U-��f[��N��	�(�H@t"�̓��	�5�ʳ�����]jy<ҡ��O_	0��������1h�T��d�30G����&��]n�������������D9r�m9�`yR毸fض`|��!H�*��?s{R4r;ήL8���꿙�4���Q�Ig�����~ׄ�m��\֓�Խ�����|�+8�~�T{�Ś�p���-{a�Wb���Ȱ���D�K��j�DNLD�e��Ɨ�������5 #k8���o$f��Pl�4%�(pC{���Z�@=�an4�!�e
6S�[o�w�9�<�C�]a��L~�n+)ǖ�F�ݵ�g瀫�,v�9�Ll\��s�.��2�S@�~�Zun�y%�uӂ.�K¶]������+�ʋ���W��L�۞M��)�oѵ!�����~��IԖ|{�Y�=�cq��W&�|$~�d�mrG�c1ChS�����`���Cq)J����3=[�^��I`wK�ڳ����נJ��AV��.A}�_ߕ�nK���R�M�s[z��.C���gs|F6�<VtK��*��2 m���i��od�>6��QG8f����\�k��g��;�DN�N�`[1� ��3��`�Z�u��>���Q6�k���_��� ����esP��p�%�A�+�b���qA�n8y;%K����� }U�I@��d5���6Ai��Pm�B� �qV�v��i�B}$pi)C��Cx��\.�R��	_�K'�ti/�B�F�YX��;7h+�b�/�;�A�Vu�fk������B#�^~Z+$GcT�&��~h\5�Y˥��;�mf��*
�i�J�FUe�#J��d+}/j�E� =nI>i@�����X�?����	�wB���p�O���ڏ�HBA1��*8t|���V�<"jy�*��W�y�➥<x��]�Ut�IՂ\�G��N؄�Ġc2��#J!�����1��"��'�7`2�h�tЖ,��/��RUñ?�7�_�w4&�l�9RI�6!��2�� ��.�����bҴ	��a����� �~NOf��>ϦR�MI�z�o���� x�>ڂh��ʄ8{�=� B$Pv��)~�r��`�:5�	l��wDs���8��}P������P;��{���):���A���N6��(3-�T�\f���P���O0k�"��>��ߍ�#��"�mo�O�ciH�Vϣ�ư��?W�~���O4��S�|���������NﭺQ�tb��J"�S���/[2�,$�>6Fv�<В?�ՠ���O��F�����~��S�������9�o��Q���)�\��}���ϛ��o�ϘTN{��¶o4�鋀ᆁ�OeKrvTԜ�����v��6|ř��,z`c'��X+kt�����%���kّ2T�!axդ�̯��]���H.;��=�����:���:U�]&G�j/��{O.*6�p�ױj}㤡�p"`{u��u��--K�W�%%���r^ަ�NShK6��=��I�n��#q(���7E�����j9-��Ei�L68���pUaj�U���/�J�G���Ry��Wn��@	Hǉ��ȧ��M�������1(���G���fz�G���G����N��5�t�����v�_[�JB���GAĊe�~�
�4�C�Y����2��Ǭ%c@��1��Bq7�y�NJ��}��[t��C?��FIQ�k�6����z�S�x����9Yh�~���J��J��䤿)�+�'93-G4T��k��Ƌ�Xcx[��{6�$���1����gp!���1����vN�|y �@�#�(RK�Q�������<i̠���-")�͋z%y�� d�?u��Pr�M.ӲO�e�/��u����ڏ��&K���^�d�)�>bx �.���C,2ն�@f\H�b��C��� ��c\�T�-�P]��������jf�6�`�T���W�5�1uHtO�q�b0b&�S:XL�E���vIKlA�[a�Z6p�졎 O� jBd�<a��	ԟ��i#��ԉ�ӂO���I���N�_����׈IL�&)�	��,è����?���r ���Vt�6�5��E[�~�V�ϙF�>R
�_|�g�h���D�EDƽA���!4�͖c��r�@[؟����*n?�r,=֝�Ze�2��GaR��&7�w��?�a���.3�YaL��!�7�m��� ��a�p��9xKKK�'`Ӛ�{�9�ܴfW�*�b1�Ϋ�f\�b��,l��"��9�c>ѥ?�{6�R��=zV�Y2\=1��_��ܥ��Z�gw3ⲯ��>���.��O���μ%Gi�zז�B��PaG������"˩1\�U���<ϥ�/"`LU/���}tG��C�cfn��b�8���PkgULM{�]���9x��^�N�[;�-�������w�XH)��ϻ8��);ɡ|������*���.�<N�{�A
��f�=e��l�b��� �T�wQ0�M5�c�|'Q0��$�p��j�3Fv`�
���*M���Nu8��������y`Ay7Q���DzNKE�8
�u'ik�@�H���3ct�IXI��:+f��
7I�>�8	��1�V4&��x]��˞p�R����L-��{��EK�A�
 r�j�VEW�%ȃ�8����%n,E����n�X*�{�1O( �	|�x�����4n$�C�=�A^����	V��A����	l����������W9B�r�EV�Z�o���t_�{Q��|.N�Z��$��|�G��έ�L�Hj�b=�*�D
I��\��$+��a@�V��wŨ�1��v7�e��_*:o�B��.���Q}皀�}Ҟ
��ڞFcwC���K�.I�
��xd?�ۮc�Ϭ6�����z&�Dfr�W6A�/@��2����㼚ʷ9\s��x�o�^ni����h������1�Y-�u�i��h#��T=7�+��@�<�--��ь�pG�9녳��øƜ�3�5��\�җQ���r��S�G�G��G����