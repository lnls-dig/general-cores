XlxV64EB    fa00    2d50����'K�պ��Eh�򓙝=��ع���W�h�mג�N�4\`��F&�R�o.�?�"��R��_>r7�ܒ3V���jfH"�ww�wa����O�_�p�^�<��s�43'c�a N�p�/oRY���%1���Zx|ņ9]Le�T48�!��Q�@,�-�z��"��G���0YlM�G��g��G���V7��Q��4�<�*{�{C���J�B]�!��xg��*kr�ٹ�R�7AD�*�f0'��<#�H\� ���!;|]$D�K����>���M���;��}�@�Č�όxF���QSH����D|s�h�5�DH��pt��Ί3�"4��G���;l:�	��B�/e~��^�!�lI�\#��$jH��H
�8Et��(� �2(V[uV�������3iW:�3�NS�η���.*�&�,������1C	f
�R��N��U�����}����km�/N�=��1��9��V�q��s����IX�_}ѱ���9�_E��-�Z����Ʃ2�v ��9_�����Y\U{�%���<�����>ʀ�Q��Ã6\a^�ns'�q˞D�V��]Yf�ғ�6��"��ƳΠ��Nf/�p(���Q��[�\P�G��'	�`����I9R`U	ޅ�_�:d����΄Ae�+�ts�r�Wsw���4�ҩ�S���n����(�1֊Ӡ@'1��cpT�U�������|^O�I��?�<dn�5Ǫ���g�}��=�/��_@|i*%�;�X1��|�4\G�vaq�9E=��3?��8�{�"��L*�#�s�	{�?�'3�c��*��.��.����:S�%��*�d~�:p �2��?���	�*-�!Do��j�n홱�[4�o���0$���Q}���̃B"�2�j���'TTE[�LY��+�}
ӵ���Q.��PJ��	pM��XO�F��;�?/��9C	rB�bX-���}�s!8���vD����b�6p����<'Dg_d ���镇fX�ҏsw�ςNw�#��n��6{�Y��!�
�ɺ�M��t�'� ����?�`��s�N�$��jI ��g�ȭ���J�V��@���i�+��E�^*��y��el�F�4��x2 �~X���lk��\$�����{��G��Ҍ���S���j�m)z�1�&ws|D)�O��u~٢k*���NI�`���������x. ��ڌ
����n�;��UD�}�{ޥ9 �+��.�9&�_�����K�� ��a�R���}�n�yh+mUZ,�������5{�J!�md� 1Q ����pU���h��c @�?�S؝�5�}�a.��Jh�I��m�-VNXh���L�o�_xyB��B Nc�S_��T��la�*����|^�|.`�� ~v6,��v~��*��9XI]�j?˥\v֏�\�EXY~D�>(��*�&10��j���Ǣ��b��C��Y�u�rw�J.6��:T�{A�^ʛ[��'����LI��$Ϋ��ۨoyj�Z���~�Ka|�R&\Dԉ�Iٜ�y�`dJ����MV�PED��\ޱ��jPڲ���R����z��0f�*]F���S8N��Qb����qޙ�*� '�~*p�=�l$�d������Q�J�h�u���(OP���$��̞Qz�1�8�Al=	G���������̓��V��B�h��rT?w!���%�1�?��Amk������)���c�.���A�m
T����'�b�ɶ��p���~����Λ�3��n2&a �.�m�et��J����7�U��uw�Q��w79)�T�.a�󣑢ޭ%�-}3'@7�WG���?`��x[�Vvو���.C�����G�f��ēZ�W�w	vn��.|*9�cV���*�@ec�]������ ��a��������~w�װr��d�ϼ���6�.@����G#3�1{�s��6��a��FMןw��뷱�CL �'G�����L�"�/E�?Kv:)6�9�����g�З�����R�$$�n�p�kd��2n��Ý�qm%j_c$�?b�>MmT��%?�9Z#��G��X��Vo^`�}ZL�/���?��k=�|�Q�
��p੕.��lR��>�?�p�Lq^WlS�1����Sro�-��Chs��Xo�P�r�[L��O�>�M�MXƥ���ƿ1s�w�Nd)_�7,�]�,1^=a[��^%��g�=��3��{�E�7�vw���^s5g�0����Z3 z�A�6?�sy=��-��7�q,��@k�d�P���8ZߧNQ^_?x���S/2����AT�#ց9���q��\��;c��F��ޤ}�,,��]y��0i�')2���fܷ .��Y�0X���{F��ut'Ar0�� ��}�����jo�f�m���;`��i���׳5dLg׈4�;�^�#[ry�m���v��`���a��QUK�.�@0`W!` ��]��:��A�rAk�Ks�@���D���l'�7Ze�LQ�M([KODJ����v�@e��v.�*���XζRX6�-�xD=�����ؒ�v�фL $�+_TU~���xb�������Z4-�q0���_i���Ǻ���+��K��|"�5&�tqc�O�Wz��.�kN���BKo;��u��m:�hC+޿>��8��Ǡ}��j��-�e0�w��~�l�(���=߃-����:_�_�5*�)�S6>]]���v�()�V+�ъ��=���,�I�Z��Vv�5��plhR���eu�Z�~e�C��m���%�wR�U;���u�ʘT�x��:��C9�Φ��t5輗��}6eW���������,�J�~+� ;�� ��t�EC{+�fG�{�=���<1�A�:4P�=є ��6�O�����O|͉�M\����7l#���>�2{/�_b7Xk�1Y*R:��P���oF���ҩT�3S��S��"�xY�D!B��ةƅB���Ȫ�3R~�~k�d�f��'@�.�v�t�)Pf����`�6�����w�{��dkQ����-t`O	0uŐJ�����S���!؅����C0r!Տ��葶Uѵ��)uv$������2���@��2_����ԤP�K�ۨ �����ط7��t�Ȓ��~Y�!B|���W ��ژߢB���yl2ez�C�����-��0�Czs�B����Y�l-��.c��Kc���S���ƕ6]@@/��#����.,k N�+�$n�NZJ�a��l[u�Wgh�o�(7n[�5?f}�ǵ(�\jlH��\M�<}��{���nc٩��ԡ�\�u\u�h�rS�� y��}��~�x�85)�,�͠�*��K��x�,��_;���sҌaG��l?���"2���d��#�{G:7._���+�����TН���9�?��p�6������OH�l��Ѯl)UC��7 ��L������Yw���U�͖�֏�C�R,�Fk�kV �@�(�?�Q-Z@Z�o�r���^�������K=�D ��� N��^�c����]N
�����c���A�k����}
��A���{���8� �o0�������-����gŕ�bI�wN��;�\*6`�V2���P <�F�)��a. $��4� �7K�[u�.�d�)�#�'�7T��տ�7�ca���J�,S�76���ӓ�!��V�9%�w)|C�jqO��z�}]Ɯ�4��͍��;uɩ:�<�t�>0̦l,���i��:s
2�5���$T�����������"��v{[�j�RGz<�����IB5U��qh�����x7b���l��V����x��d������Y汊^�؊rQ�z!Y�Q�3.n����H�?�. ��*D�w.6R�5gl �F,�������X��y=��:��f
��b�r�����u�櫱�D�	�8��J^X��B���%��8=��Ay�ʎ������6]�D�g�=��i��C4�2���[���<_�~�/r3�_���NnPW|̢�b��Q�%�������d��s�.!���?�Q�\��� �SҘ�-��!mr����Ug���PnL0fAk�����A���qEu��j�J���w�V�cɹh�@�_Ϋc�*e�X�;�x��<k�f�9ꮠ�h��:U=0��"7�2~!5�=�{r[pR�33�;b�{��B3B�D�r�$���Q��s���@(��:M4���(rϯ0Ⱥ��f��.�Y��+�"��[x��f�}G%)y`��� �P��.�Q��B���┛� i�O�R ��c0�Hf�1���Q�����U�����b=`��(P/�Z�t��6�Q�0.�^�3�d��SR�V�����hu`M�lT�|<��S�N2�j��%���xa}do+��{MhDr
^澿�P?^�4���=������Ч�tMeJ�d/�A��Rc=q�)6fsh'�@�͢��2��*��`��S�VCI�	�F����12�����;o>�
�.Q�B���
�(�4ޤM�뚉sz�@P�sR`��Ku��O[&q�J��2����1ȵƖV�
��lS�wI?�(bE�N��uK��u�#>h��0��L'�~|���q%�r�J��'$|��T�C>n��5��9~�Eu*k�6���˧V7g���jLET�[d *�H�b�O�H�~1��5�e�!	Uc#����5�^�պ��)����F�`�3��[&��Hp�F'��j����گ�ߟ�Q��Մt��_u����YjE�o@�X+R4�N�V��j�~ҙ ����N�{����)�c9�e�ew��jc�l4Yظ���Z�3��M�u+���s\?!�$y�-0���wv�x�}�
0`Q�F����Q���믷������I�lG���k�|��*f���k�#�J*��U8�g�����%��q �#}�R��l�׳��P�U����R����'P�b�E���;�.x�̀hK^U'��	��Bi�K�Z��Gi4���MhǙ^L���'`󍣕嚶�j��~$ٵ�2�.f���Ԥ�`*G��Ȉf��)3���xB�}{z���#0h`��Y��j��֥Բ<�b��YE�~� "�������+&���=�09���LrYu��q��d��~)4Ҥ?`�*����t-F�B�w�>���0Ch�2����!O^|��qF����䐩�Q�i��n���$�-�4f�����[���5�<�u�f�b�
.�8H�׭g��9�ʧ����7W����F�ȃN�U�.�q��ϰ|�D��ՇB�|�C�"�x���ޔRLS��O>�Pb���L�hA��]�`�ͮ��&:?-�P`�w�w|�xo�2���`R|�-^���n��C3;8�G�3�jI�� �� ���T���<Z����Z��F<Z {͞��H~sL'9�jr%��BTL��@o�)=ͻ�Q�`}��H�?�"�$��f�zTL?�.IH����F�8�7�a ntW��f�H"�}�-�3|�c$�n��f^P�'��I71��q�V���e��k��6� R5�d�r�TucA��u�-96��Dd|�І���阫z]nBr�YI�Ke���p�y���Bh��S�p���o�ͦ�;�࣌���~��o�p���Z{�#~w��o�)�D��l�&Hu���ރ�n�ڃ��'%��`� tD��N0�6����Mԣ���=��������Y>0�;��J1��L��<[+��dr}��O��B��"S(��jfw{��.[f���Dd���U�}��щ���k�B��O��X,ק��V�8
�C��@���
 ����1�q����Q���:C��0"��+Ԡɿ��z�҄�z��hK�p)L�����k>@�\Qo�U�٠s�zX�|]�)�Gb�( 4hJMɫχ��T�G']��O�?����=Cș#&Z>�/T���$T�n
���� �j��A�s�%B1�V�L+v=��KqQ%X��ic��xo?������(R8mi�u�%��B=jUs:[�p
��Ñw(�V����@ BG����%z�+��"�1�cnW�-�DS��K$@80|p�Rp�[��g^]�l�aQO5�3V~����+�,F��<�< �̪u�5aݶNC�C?⌳�ޛS-o���<� ��[�4���q,��.UVC��	��7�5;�!�s>�N��T�+��)�RG2��;}���AƏ����	����YMv��🿊5�,�¶�W!Av���׋f���J���#�u/�K�M�Jw�A{a�k��H��D ���AHLՏ��X��)/5�ş��������	��.3}�r�_�=��)6�����j�����֕���!F�'��v���S�t�(�_��� �#�^;���EԸ�֮�;����c����p�mX4�}5L=��1�I�̼-��&��� WD��G߬΃ ��f"��ɄI�V�h@0�eb�z�E�[�d/�֢h�����@�&~��_�S�3��pt��~��f�y|�u�x`�8�񆵇�n�|Wt�U>��Ֆ����~�C�(�F_�����X��U��)���	�$�<f��D[���~�wg_��<�?^�4��6��(�������.*�*�#[@7_f�h����!_�,O�HK�Z��ڳ�5�)�@`�og w��0lbu�a��u��h	Q``A�>����@�dB,J������!m�kl������D34,m�GYo�l�M�%�-HY�������
]�W�py�Z�߭�>ySJ�W���A�[���2l�-��S�lI�9�~}��`~0k��{U�ܞpT��oFQ��Y ?�����hw�� �Mw�MT�}��
�d%����!M�T�y�޼�l�ejc.�罃椢�)��9\�,��~`�'�@�y��BX_���k*�`��bc��@-�]��ۼb����!��|p�)NbCo�z�{��M���Z���X�p�?^7�J$�+��j{P�w�~G�
���`K��h�1���*&��1�M�!م������j��K6@*�n��Ձn�ج9WA�'D�b^ܟ;a�E���B��-EJ����MF){R3.�W��C���:>�"�ꠏ�e�B�8����"#�P�Ε�k2� �֟J��M	$@Πۿ@�l{���CJ��:�.:A=�ox�������f���e�3�])#\xa�+"�	���L�b�7�,L`4�5ݓy���0�A�v����b.��P�w���2�{�H�۟�	��<�U��h/��?�1TB�	Wq�*�lc������#�<�ڀ��0���n6����W\�"�`D��� QJ)[��R�7���
ؗÄ"�v`�5u��?��Oxf+aI)���HC�șZ�&Zߡ����&+��{�G(��U���a����re\q�s4\���lX�!-�%�>/{E���T��:,�|�l�Xl��ϮGc�󸛘������x[� *������lb��h:}�0·M�^±�a>�Q�',�Nе���Ue��7ҢZK
S0W�k{U	F ��V�!��/�}���|�]�	���:�����#-h��\�ܰS��P:��񇜱@eR�'�^���}�A�u�W����ƪv��,���m��W�+����F.S�pL՘��^
'��lx�-�U����=)AL,@�9�"����U�F�UD�o�m�W�47��`
~�3*��_L��A��b*���F��*�u�5�	��jV�*v���R�r������E(�����-d�=<�Mf�&u�?[u��������F�ݧg��|�Tv���R�ܨ���Ѻ����k�tЁ�skȻW�BYx3�3�%�0�k��Gt�ͼs�Ode�[U�+!�Kx���k�\F�����R����)W`��%�{ˮG I��꼟�k ��8�0Q����Ȳ�m݋H�<��(׶+pB�B�O�tl�z��!���>%p@#�[�p�T���%���B����C���)Ԙ^H�ě�������V�Υ�K����B�LIOT��K����AȲ�:�{A�gٍD���w�U��ɚ����iq���*f,*��i�q��:�,��1��p-�k)Z�4��d�{�@�r�sUsa��hA���r��W�������L���إ�>=ز\�O�dV@�ɩ���~�4�.Z� �ЙllJ���ڮ:���oR�Ǩ���ü��v��i�n�et���j�p����~E@@����_
˜\�XC�X�`?�p�r���yX��h���;�)@�U��y���_�.a �- ��*zyN��V/r�����r�օOFW�������$N���M��{wF�S[Q��u�1v�Y; ���5oM8+XY��}�%��4��ł��/<1�V�%�g�i����r8"SpY�T	�s2�P_���W����h��~	�45��>�]��2mځ�n�Ou5̞��P�٬oD{���y'���cq}]1uAr�ɢW����T0���Fs�Q�E�K�K�j^��`�u��9��#B/�l�Ԑ@J!�T�/)��A�8��>Y���I���%vy�[���;1*�8�F���Ft�zW>������ub�m�e�a���uQ�
d�Ay?�
Q����I�{�3Xd�d��e���>[ 0Z�t|����5q1��LN�R���c��#0T���L���+ҭ:ug�vd0����)��#c�2��р�K�F�C�L�����Kn�����v�5?�F���X��\�QVq �]�(b�o�!�SN��ډ݆�Ax�e=t���4�4��BSɺ�uәX�Zs�i�H�4Zu��<3Y`D��Rd�4���I��9�|�X����tg[��棷��:�+���(�=�,>�K�;�]�y� \�YXb1��{*C�	����~n|yN�w��h��������7(�_3�q4Z4��ܿ7K�x�p��z|�⛐s>�a��2��>5����잲���G�J�n����0Q��ցx\�̟7�{�w���仙�}`���f��Dl�:k,�;% �}��gj�E]zy�k��.'d|���"���?A��ۑ�����eS���0`7@G�nZ&���g�a2�-��(ߣ.���^���ZS���U��{s�-�; �`DhX��i���������/RL�X�[bN�^���sH�W0��������9�����SY�Y�r�/X$YuUZ9�5��U���b@�ZO@0��*k�J��塞� ���Wc�6����R�������lKr]m��f�NTG�y
Ò��k�r�E%h#��/�n$��v�o�g�z�KC֫(��:�4bܯ9V�X�����cr?��K]�s�{�e5V؂Q��K
!�`z�~w/���>qL�i�X�%.��3��������  J�|�Q��0��O�#��	FI��	l�x&bWXH�Xo�I��c���c��T_U���fåN�L��Edʻ	�(��Է��R�26�ضw�.��@@fK�w��x^�o�������0�+��a��-�@c���[�t�ܵ�y���^o���*�ץ_E��[�V���5�iu���3%�̵<�xu�~����jM�]B�ʓe�D�=u���Ca4]��<�E��9	���0k�I�M��kn���+އI���2�~^�}�XF�*di�L-��wP҆h�W��9��R%�cE)���G�Z:�]�s�܃�y�.�p�<�` ����ܿb��:msP�5g\S[����܁�f��2>�4�`9��J��F�7�T�2�f��K��*�(����;ԵIgKvWj�e�G[t�1�2�<%VF��Ώ�Ih>!����紱��i�5UH_b��gmU�OШ�'��f�9��Ҡc�+pq��E����F5�E�_�ͣSтI'�1�/|��!�X��q2�y��4p@(S��<qz�aQǮo��lԴ�yė����('���ӻY+2<P��0"�Ǒ)��hrH��j�MU*Q[������n�Nϐ�_Ϡ�Pn��<m��������gT���g$��>������y5p)NB�zg1�ʃX�̋l8�1.�c-���;��Y4�a߯�5�彦p��{��⡯�0$����F�0ݵ�*�ԬFKs�wx�������aS{0��Z*ź��Sd���-E����v��_�y�c�qd%�w���>�dr���؁u�����'-�h�j�eF�p�02�E�������Qk:>��F���>	�
r����L9�^��X��L��H�n��q�h-�T%@Y!�����M�GlY�xmiz���������im�R'pObq���G�U:	�&z�o��[n�W,%�I>iy��x�P��<��� :�R Pp��Zh�����8�{��.�D�a@"�᧳E��@^����>2<����6�U�j����
�Z�w�KL4�n��**�@�^�6ն���-�h͕Tx>!\(H��:�p�s�Sk<�_X���ѵ��&�gw�m~T�l_(�����nIMk����ڽ3���������8�`�^4��22'���kMNN�*{�շ\�8����W{@���H���\��x����֢ _T�c4�k��9����p��G����D_�2ү��h�}\�a�-�MuO�YNL����R�4"�"41
�M�
��H�n[9���n��*4��.a���jd�G���T�4)��%��x?љ�8�'���/gG���B��B�U���7�A�"¿Sєx���O�.�;	j)˭�^�-��Zr�p=�^�P�亦��~	��I�h�v4��۽��7�D�+hF�^��!j���P�;i����D>��"�a�&��{_r�)=����cRg%�Y|*�93U5UUn3 ���:�m�|nɴ:����Ы��C�w�E������#n��c�z��5zݭa~��x�U�2>�W��c��^d��Y<������综.��M�.?G p�VN������@���S�M.C��Gm�jt��Pyp�+����9������x����ł8O�q��.
�+˔E>���d���H��27a�`��}�+Xw�V�.
F��B�L��'H�7o��[P��a��Rl"��^p>D��M�#�@�Eֳ���V/4i-�a�g�s"�@�9Ct�6�'G�S��Y�G��]�i��-L_Z��e%���h��ޛZ��&5#�b������i���QNXZ��ղ���et0�?�Q����uL�؞��Ƕ�7���1�������:=ف�#}[e��[�o��q�5�Q��_��=�d9��Y"�������s'�Z�~�MZ������m�7�@�>Y�-K'�85f�ŸP�@��FH�.�Uٔ�q$�6腖�[pĦrvy���Q�(�u<��S���ۥ(�g2e�
8v��_���=qͮ�u�4�9v�u4"������� $���*�ѐ�XlxV64EB    6552    1140�c�3-�h���18l7�ɧ�f��5��㇣��]C;FhC�K�el�� �����]�iD�W�A|Ad��\Y�V��a���^LA��h��ΆV�p����P��=b:,�h2����=98�.?�G��R\ei-ɚ���k��g��[.�]�}Q+� �E7c��2�{��w����@!�I.��P_������*��ƣ�E�Hzn���yǽ�z��х�Od�����Fz"�q64���	��2���|6T/����W�χ�\�.$d�K�Kn���l�~�R���H��fH��&Z�'�.�T�>EU�Q�*i+��M�zIqp����HС�-ŋ��������zI��9|�w�C*��t�+�gc���2P/3/Q����� ��r��ZƷ�;6.Ձ��=�٤��]1 Vp��д"*�x­[�s�:(.Z*�Y"�+�m����#��h�1B0^���c��'x���C2l���.�Ɠr�o�&G#3�s��˄:���ε�:%���ac[l��\=eGC�Ɯ�X�5wK�!28�5*qlT�_A �n��Ha���X�H��;��:}���n�!��J�7��q�W��K2-����]aO7{�7��l�2Io�6��ZPv�+L�L�L������c`�}(�zk.���v$��$�Ҋf�b8w�v�&�6��/�M�
�˴�F�n���}�X&*}1c�Z�;WA`y�;�?;��r��Q�*��y�֕����)��ZW�/�d�G���\t�;B�n��9f6/-�uג�ff�2A��\�%�oI?�v��=���_	Q�����ͯ#v������_N�==�����p�wF�\����]�Ag�LO�/�(Q���"���\��2�d"�H:Ɋ�u%*���S
@J�z�	<k�Q��^j�mр��-䍪�O^'�NyV.�I.��-��.)n�k{�:!�4�Qq�#2��RʑL>u� Gr��7D�_)Q'�Iƚ��,�:�H�v��s�nE��b��*G��,^e�˛���U_�c�MBx�pѤ_H�*�]}3{f{��p����H��c�,�@��(�E<��t�Y�py^@`�G�]:�2�-���Lt�:B?�����k�r�c���ˈt(�� u�*����������@��w�4(5:����]�(.��D����ɈЪi�[Z�oK�E:T��>�S�(���	��ɣ���Z�
3:�z�[�<�!�'O�@�pȢ F|N��=�A`�~vV���oMı��S()��f�Ө�H甹�<K\��ϼV?��Ƹ��8����=���ߚ��ѨR*��쑷�46��|�)u��G*5���9Um����$������5�Q�7B|B\��^�O&8��7��X(���k߮e����\���\�
$�	܊Yqi?����;�wr��D����+'��(��F4P�䌝a���?^|���қ���,�S�*�Zag?X��@)7����$��W���P�Whz�l���q��Mde(��f">����$r27�}��j�4+��d+�t�pf b�`J��t��.;��u`:<N8��J)%ҍE/k��\�&������ �?�_Ƴ��ϲ�X	]���g�둳)cę�������0�����[��
k�M[�pGh���df3)��k�[@v�Ho������HS�:E]��{%ŦMl�;̜���F�7��tJ;9>�+�¬D���Rp�*\�;h1G�!���[O�	?�����EWг!c[P��h�0�9��3<h@ �j��<�#:䖆{;�V:�1�E���;D�(�o¸ZH���F����E��(s�ѥ�
��]٨Jdq�kB�@��H�p(3�s`�3;�C�SC����nq�	e�#�)��f�o�ϗͶ�O�f/d������,?�� ,1�ǋG��Ϻ�'`�aa�}��Hǅ�#�7?M���P荛>����>���t`�d+����p��f	<hh2�/��:iC���n��k��TZ�U&����~�y�%hXqc�W��	�gR$��=��G.�8l�̓�Ӂ0����{�D̿H4?�f��9a;��X�5�S�o��Y�Z΄��S;ַFl	t���H(G�_}�\u�x���
��Z�!��|R\�i����X�h*�2�y�wOM�-�2�̂�H��;�N�1w�b,��>��~��k �������ug9W�x��$�ܔڏ����N�������*�����q>l���~�l��ZN��`k2ᜇ%:ϴ�Ku��N3�k/E;=�:6���<�0����;�?���&G���l�����"d�@�u�2(4Z����c��_{�]	�C��@EqY[�@ɍu�_
&����?i��������l}ͮ&��I���T`G��]�����ҡ�����`�4�pF���h�$�����[y��㶔u�S�Eī�^�5�@e�e��[����/ɖˌ�^�b�)?ɞ��1�!$�#"͋ÚP:�A�u�7IEn#6��Œ'���:�I/�WV��_�*>LH� �!:�tS֬��T��%{s���E���W7Ѿ�jgx�z�}�%�?4.�o�F�FW���Hg�u��V :C��	�93~�Q�!r�X'�cq�n���C`�qSЃ���%dp�+�Ի]$M�!����G;�p�z]���cw�^ �"�pr
��w�CVG�E���	�}0�\f��K���u\���ެft��l��d8���ja����O��[ZE�j�;)�ϧ��c|����ҀրƉOe�L�hZ+�\pg�=��{�i������MꙟG5H'��}t�<��j���6����Pݔ4�#ȍ0��5̅�cx�t�����\�k,r�q�i��SH���c�[wB�v�/RF%R?�2��t�>R���j�4X�m�"�;��i�q�k°9����fM߃����A|I��u�-<�`7�	c~���<(�+��Ґ辘�y�r�G�S��f���)0�Q�N)�����؊���K�8!JL�B���K?�Y��I��H�fm��(���tо�O5G���WF�C=����r������6��x�)b�j��#7�4S/b�P��w���j����@��3�ȁfuda��Tݠ]H.�ϖ� ��%���9K�9���C��T��n����&m���A��U�S�����c`������	I[a��>5�`\����4~�dC�Κ �D�&S��eB�/����Y�=&�&7E�<�˷�i1g��X=<Y�&���YW�)�+(q��g��h�#kBO���ۣ�r�9\��' :gR�4]K��r�0#��Z�hr(�z=z�<��tg�=�SS~8��~��`��Hj���x��}u$��� ��W�����QB�:�ɟ/,�KR<��Qyb�Nq��hnU��|�8sD_Y~��0�% �wC��w�S6�����|C��|-�`�)D�cЕ�ws�m��L\�x�Μ>�3�o?�V��ͦbM�G�P�������g�e��.��}����)�4�J���K���w�P��2 ����8�M��r�Į���'~SQ��-���ϴ��d2UT����z�Le��">�)�1`wf\�qUP.�2��?�F����\���j:d�%E�0�#-J-C����X�we}k�LȎ��.S�]�+���sݠ��}T�/VU����?�`�,�"['�L���|$a΋�����+yw;�gY��m�i�DP�ʥr��F/o��Q��� �����OP�mt�-�e�J�wd}f�۸~ȶ6���psw��EqBEI�I���Ŕ��V莛QTfD eqnv�\54\s����a�	�voe�U��8�ʛ����_?�۫���%$�S���E�7��téG�f8��<J�h4$���΢���u���| �BCȗ5Gΰa��a&懈��_݌���r-:Ys��q�O�fcĦ�iʓ�/�dj���>���v�b�c��û ��VN����v�N��y�����j�L�����6�lsy�P=
A�1sI��H��5�n���	-��Ek��4��_CW��_�v@��(HK�C�<�^y�ZS�+���׊M�ۦ,x�ir�(�Ӿ6cH����j{8r�M�9�r�	ڈ0vr�&�x����-���@��f
3 V��
��
lCrΑ��Jd���r�t�~eg8�ǕLZ��G�`����1��s&
t��]7�uUM�����$��@�[j���$�*5̔��wس�*�\��9Æ�UY��Ae�{�v��:�oK�|	\�Ы���G��8MUh�L}���)RP�����Փ!'c