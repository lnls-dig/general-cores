XlxV64EB    27f1     af0�@��Dek��'hX+Q@����gZ�G�҇>x���ǀP�<X���|o���^���r���	vz�졩_�Q�(~/�=t:�B���(mE�D,�i�ط�qo>/�Z樍�ؿ�LO�«�#���+3y~b�X�9i��|'ll˾��%y9'G��};x�q1>�*��_c}�O�O�������f����3����oP6��t~?fe�C/�>̲����qS}����<��x`$.}w1��{��h!�ϣ6-�����ڻC\��o�!S��y]�
�Mt�'& �5��RI����="�P�K��$X�O����wZ&2B�Ȑ����>XfEL\.�;Y���rײCҪ�!�-�t�pҪ�a��
	���Bs���N1����6Y�s���Q/
��_Hz��DY�Z�B�QS)X��#��t�x�uv�<#��ܢ�tc.��'7�]#a��Z�F�u)m�m�����k���X`k����$G�����JQ$-��ǃ��0o	͇�M��.5�Z95����� �L��1C��*)��Dy�1v�Q�/����H+�J�{b>?p�x�!!F ~nsh%�ܺ��<����oʾ}6*�F-��m�f�-�w~�(���ͪ�S��'�n|�����Ek����$����' �aA�mKͬ�(x
K�YE.���#�m�B��bF��7��ǹ;���G�/�>@��!�7�'ȓ��d������61m��3�`�.V~pL���:��$���|#�	n�� 
6qS'�ȹO���J^��j/��sW���m���*���b9�
�~�Ԣd��o��P�Ro|��e���a��{Zt�NUv�)])<L�`ÿ�&�D_<�w�q]Q���ɜ�&ͷ���<�!h�:C�Z�� ?sOGi���^3�e�"�K��	=V ����ߴ`�5����%��7�?n�� ���e3�t�QMy�n��g�����7����.��9i����T�ջ!/���S�����,;��W�ө>$c���zW+\)+���+�X���^�:���g�ԖU1��*7u7�аp�&��P����c�y͊����Ɛ�M<���f��Ά�?�G�U�v�#�a�}�b�5�帽��*����ӄ�6�>�wY��:��{�%���-t�e�U̪��'�{7��J�B�Ֆ����HQr�*���I�_�LS8����K ��s��yū�������� ZDN�֞����^�y"7�W��~-i����粚�Nb�o7Y�4�T�mI�mu4���0B�C��T���hRؾ97�!��_�|6�	�QvA�'[���H�'����2ylw�.�ɜn���؄���w@�������0y�S��xA��"�=�;`�J�x�C�`�^���>Ȗv�a�ǝ.#�1W6�k�z}������i�D����k�P�t�8.N�i��fMD�\ye���h�o�v<XJ�x,YN�q����N�Ԣ6��@�p�}�$}�J���B�` i3����㮖Dr���æ�����ڀ����;%Q1O;Y���W���4@6i��O�]�O})�� ���:l�����zTn@�x��B�����z��/r����FoH�Bۥ`��o��aN&����g�6k�С1ܸb'��������ʞ�b�[SO�_a]�xx��&аM�&��us�@����N�=�?�(#p�+"8JD�Y`�
�]ն���j���E�K[�v���;��hbj�l/������)�9���o�"�w?�X��I�|���
<Sh+u��,�����I`���e
��0�9�Rm�{��m�딸V{S����)p����Ƹ�'�|6�L��l$p�Q�u��GG��J���'Z��I�AWN3c֞q>@�^�*�Zk���e�гg�){Q.ॕ���jA-4S��n��iu����~�3��~	�.4I�ܘ��v\��y.����9[�"a1q#eC*�@D|��F���'�E.�dM8jp��+a�^�Lj������	4�(� �y�q�8o�o���S![���&Z5K�k[�uG"�{��F/Ma���p���¼���"f�5��O�����%}]�c�$%Μ/��`X��:�|�T���s*�0�M�d�u[T��նy狽�G� �*P�}E$s�����Wy��g������ J&H�v�J�-�QQ��6��"�s�0��>}��%��Vk�H����X~���j�+;H�C[AιTZ�>^۬Y��,���Q��Ӊ��W�Mo�NNW��sE�&4+W5��|��w�TgO1D�g^�8.�tHWN���IuT��9�w7�f�^�?�=j7�P|�p�(!����S �@�O 7�������O69��j/Dy/��w�)%�׀"�J��|�Ϟ^��XAjU7*�E@k����2�\�b �����$�劙��P������'���׬_ B�b��Ȋf�����VC�6(j ����.��ר�l�3�ؐ2Z���;���ٸ��R$�F��3�jDK�1���j�ZF�d
���ƿؙ���ޞ:�����,������9�]*|$�Îi�n�e�ƀ㡡~@��Ʌ���p**3�nv��lxkpv�'m��M8�?��sk��e�	����!M�t�n54똲��U5�)�������K��������"�ž�2�|K�ݜW��dAQ��wv�� ��C���`Zc�<1_��0���J��K�$����7TV;����<_��)��