XlxV64EB    2cdf     b40��?=y����T5�����d�GH*h��x�������9�.v��_308��<+�Z9��E�Ve��'[oh�.��{`��	fM��T���,��
;�Gz�Y�;��		{��T�u'b��C���?@��*� U8V<~f�����]��e�+����8 n���ѯ<��'>���D��诋sh�Zx�#Tu�o,V��PXy'V,D�$��HZ������x_/�O�H�X ��VU#�Ǩ���y�]�& �&��7�(�wk��Yh��� }�M��eD$M�&T�9,)��nw	>O?�lu��|3����1��f�=P׺e�
W���O�Ιt��Ӆ5�W�,�E�j,"�@�kx���>A4�Vg��MEs��Ygٶ����1��g���bC����6�������p�ir��DH؋��@Oa��~� Tz�SH���ܯ�����}���A�j~ms[�"�G$�_r���c1�*�{>�ysJ����A�{@�|�I&��!�~J�F�ޖm�Ā��	����^kͪK��7�}�DANBjaߪ��*��T��Aٲ�z:A|�	źA����$���;ɉ(;�?~�='�w+�Ra�t�V�����0��������� ��=T�&�Ty�~�V7FT�&J� {��jo���_�uM5Dr�7�q�����M�d�>r�m�u��0����ct���	 �1�Dc��=�F��פ'x�Y���V�:V����� �j���u������(N�l�HeF�*Wx��pl�)�I�J7j�j���=v�ì�d��7͗鸎Ӌa�����s�5i1����kY���w�Zh���e'�P��S�+ѹ�M=�[�z�g�)�����qC��i�5x7fd�n�몦r�яi�cJ�SΪD&>nAT'qeV���|��Ht�P�,� X���P��:!�lD�ao2�	���+�ֱ���Ro�SR�3��sl��^ ޠ��"��Q1]ls\,�o1q���D���KJ{:D�ˌD9��g�dღa^��ü�Ǟl�`��*�!X���wN�+M l]��j�D������ZgصUgd:h:��oJ�����b��D�&���sޛL�ܡ�XzX{9��X?d�i!�k��>�(�zI�/���{{��U������[�.㌍��rN�*�=ѹ�b�L5WN˶N��"AL>��-���b2x�M�®�M�m�)ӗ'�Uhj�!���;��ۤ|��")���Rf����k��m+<%	����J����?֣��%���Lɑ[�T��CR��G�	���:�d�&��?�r��L�Ä�����/=&�Y��ɱ�@
s~ �۳�&.�ť���͎��X��{CW��)�NS�h�@�I�6bR�a]_��haUx��k���X�����:\:Dv��Ǭ1�/_I���4�c1��@��r��;�c8:)���)��%I\"F�	���Z_�s?#�Ф���Qӏ�U�=�&U�"X|�Qw��n_��$�9ͦbv��ՉA��lsiG��o��N���C��3�� 6�*c�&\Y`�C�Ԝ�7
�1Yz �(�/R�ꬕ�F����!��Ɨd+(���I��������$����B�Hl�w}�s�z�ȍ��UY&VW��e���K�u� ��@�˹���O��!����|žZ�������K&Sw|>O�.N�(�V�o��:$4\Z�����P:�s��e9�	1lJ��-��3,�������=,�vs^E�!�)7�**JP$TN��=�����H$�il�bS8������i�^/���}K��yUu�tc�u����%C�{_�}���F��Z����6��r��(�X�F9!)��G�Xr{q%G�����@Z���7�v�[]��l���]��p1��PE����L�qt�V����3U]�X���B��]�OGjQ��] ��*�gƹ�T�ZӨ�ұnP[M0�(�V�txg�E�ui���n��xU��g�78��n(U�� Ș����(�[�1���E�u�����|�&�&�!b��^��5=���#<F�A��}���8�N�}kG�������_�b廔�d�<�B�dO7.�m���kC�ĸ��zM�ILcG����#좀	�m�x���δi���hE����V-WP���Q2?䎨��5͏tD�����cd.��	cI���&bt?<�"I��yK0w	;M��2};��1�^�'�-�>M��r�k�$Qb��u"�1�5yde߿\��f� �7�z�{i\���C�!�"���#���44%��~q�����kë�p:�`��9�c`�U͸Y_���+���`(H�;vMIф6�<2�Ρ�X�I#M�%��\�x���B�=��I}3��B5z�(q�P�Z� �N9��ߔ֥F�,�ɺ{�}�PX�N�)��"��e#zR&��ە�����q���=�r�.'a��,������52�-X�&��e�E�@�Nd����+���N�A}�׭��8u^M^���	���ɔ� ]�� ��P�M.�����G��]1�S����"��}��/$?D%����e�qļ�2����.����*��T\K�Ӭ�uz�/������ BkKK�T�H����M�M�(�����ZD���O���:Hs���:8�LcZ2.ǺL��+��"������6�i�����g�g�mL%�^��;�|T�J\=Y-��1��y���JeȺ]�67�P�-7���@��*�F��헭�Z���T��u�jѴK[�u�cx�l��b,V��M�Eɭg/�W���M�N�W���Rda~���Zߕ����<�IO�D}�`����2��