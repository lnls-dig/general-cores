XlxV64EB    3d81     da0<����"#�(q��U��j:[��U}Ř�̡�,�se�J�=f�e�-@�J�����p�g�[n�|��<jO��K��n �Ml�	>��-A�Ja��*���֡�F�՜��x�	�n�w:�N���{ۚ�U�g�ҥ��|�)�e;A`��S��S45V06'� ;"�;�Q����K>p��H��O�@>k}���:K�� q�"n���~��n�P"��.Y����H���R\�+�BU
�X?���qS��#�@!\\n���|M�Yh�*�����oSW�i³������W]2�w8�7m��۩���U�i�y��c�R
a�BIX���@�nb��R�_�ܑLy@�wCc�����~�t����\�iD��g�����k�����Y^(w-�1j�1Oq�_YBj����!$���lC:����!����� �nF��5f�N��j�ױŜ�4xb�q�Vd�y�����җ}�XjKi�s��;_5���T\[oo�"�dFK��L儿�O(�EU�m��%'k�b�`����~K���1�>�1OشP�� �:B�^Z㢶9"f�,&���zV���k�L�g2m$F�Q�.�%�(33VV�����ʵ�.���f��u�Yǿ��$���Ӟ�3eS�v��D�ISa�A`C�AqM3�m�Ӣ�N,��u��*	�}�1|0Q��LbȆ�MA�W��f�>G�I����=�]��'P�iY�?��Mh��c{�#�;=k~�#GE�NH�P��q7[ ̭���F�:K�j�wف����HT�����M���G������Kjm�T�1�����=�+�/'��v��v����ׄ�OM���n0M�<�-)��ʬ-��#����{�b�:��e��!H�9r�Qތ�,�߯�v6<���[�S�0׮$C�!sg�Աl��e�r���7�u?I�ʋGy	(:�M@%n���F��Z�ފ��W_n�]:o"Ӣ&��}L�8~�}����a����Jy+L��c��z��Bk��[l@O��q���o���I��Z٘,���UEH�ٓ�z��6����DO�Z��$�ȅzO)��T�D�����I)I��aJ�+&��yc]��ÃN�k����PW֌�W(5*S��������7�(�
���I��'_Sqƌ@
��ۓT]���38��k�i�e^c��䥀��C��nk�);��Cg��j�+UX��9W�����dQ�u��:f����B#�+l�m�(<�z�X�#�{xTY8�m��c%G����>9pi�F*_��:���}�m4ǬM����*�/�z����\��j�՛�\�s�k��6>�1Bt+��#ߍT�$��eT��aV��x|ÿ �����#_��;�A,����o���O��~����=:�9oU�1�3yB����^E�QÓ��K=����p�,׵����Z���ߖ��؊��ݷ`b=�"5 ��ָ}����D��L ��~�T�H��@n�!Ռ0`x����g����y�SP&�`Zj�|�v�}��Ǹ���Jy;�ͧtG�������*ƺ��ڸ}B�
�S3��+�j[���#�v�7�;Q �:��yp�q�t�u>2�2�i)̴_�����x�t��O�������ѲD��S?�S͋F���^��Ѻ۠��U�+}��kY��� B�X���a[����2+��{ v#BS%&�X�;���2u!��������y�9E��'A�K�=&�ͬ���\:�D@2jD�fD ���J���dYx�7��B�!A;��_KO᳢�u��{ 5w��|=*n]�}Ҳi�{��$���z�i".��K��>,S�	.�V�*$	e�.�y��r�aB!)Bf�8�8��e>�Mh���+�$m/�gd�!�U{���	��n�>�K����+
O7�(��]�V�Y:0���/���q��Vȃ�˝H,�bT��ѝ��O�j*v�3RY/�@%|�����U[H�l�
���)�P��H�Ԯ��B��̌�mo]Y˂)�Ӵ�8���C��Ŕ�G������<�U�i]�;OFa��YB9��͕��P,��s�u��OwI����e|�r����o�P�&�M�M��6���]ȍ��ξ+���[C�)N���5���E��ײ����9h�\C��GS]�IDg���U�8�
Yq��]r���������I�{j��IP��6�լ��� ��h���='�����ż/����el�A���@��B�w���L������iKh~R�(�ӳjP@_Aml_4��ӳC�<��=��1�WO��U��8�d@�@�Rba�#��-k��楃ɍy�����n���VZ�-n��������a첳FNTL{�R�Z��hk@E�F�P9�>
�I�YT)�2�Q1�`����zP��@����.��8Wh�N]�,�7,a��{���1 ��C�LdDԍ_�Jd�N�s��}��E�o|̓V�E	�Q�cq��,�������SJ,��i'ԯI� ^�%�b�Y
�*��G|_iSjiH���T9�"�HQg�G�PYBP�}Z��}^�Jb�'[�u��L"k�2��mL�cX1���p�wm7f|j/��y'��!�ݷ��
�j��I7�yE�e�	)!�,�j5���]�K�	Ix�]}f\/#˅���3�m��Y�C�x�83�	���S�=����ވ�湃�y�A��CiK����V��R�#H�juR�Yz���鼏*�;5'� ��D�"�遝$(*On�Q�慇5VG��[θ$=3�H�mG&D���c1c֌O��
����g��ȥFB�N��h(l@�n�ez=�u�b� Y�=��;&'�p�|wa�j�xI�ym��+�h��CX�,/}�KcX+�Z�9ў�Wl?��J�#���x:n��2�w�A&������*-��pn�� ۧ���:j�$�4MAp�/k�nnp�\���T^�E��*K�S����?�Cݘ��b��<������i�3�����{CUR[��q��g@_���_n�/��?��0�x��8�BR�r$Ň��#lc�]ᓃ��[�Cqׂ�[����-� �t\`�nBY���Wvq�7��CC��oׂ�΃ç�J��b�hZ�A�ȳ�������ʨ�@ه����n6�,��l}`�>6����8?z���7>2�ش����No&NH�M���=���H��D>�8m�B�s��dLz������n��Z�j�+�S����߂m긛}�E�B�!��b�0h�Z6^8�73��{>%���,�N������ڑ���"Y-F��~�&�S�<o�x(���z��q��D�ݟ"�vϛ�N� [�� I��wd�o���`1%E���Se�n�����3������L�;	%�0����];(�v�*�ᾷY�.�g��#�����]��.��n�;�n.�8ӟ��Ħ,��A�H_Qk���n�&�