XlxV64EB    a423    1d20\6n�ZH�%q~=ރF�@8Y�b��i���̷�а}#@T��Nڿ�ҘM0*��y��C���z8�NkQ#_ �K�t7�������(A�>�0o1S����|Y�R�G���)����o�a� KQs[�t�Ueq��z���>-��o�b�W`�cRo<�����'g���������J����F�����h~���U��.9�
G0gc��ߕM���W�SJ�hE��������Y_�潸�Ѻ�L	o`��� �G`>�ҽBԀ�]zbZ4ۺbz�lU;@�x^����&3�6G.�`Q?�g�D����APx�gbsk`�~$*ٷ���|��ڳD��'
�����9>����<��&*�z<",,$�H o���J;���'e���a�&�����*��9սڭ,��H=a.�Z�n@<��J�^�+)��;��{�;p�+����U4c�:<-�g��(�����¼<)ʙ��;q~�u FG6�����@'i4�l�`�c�tM��� [�f�Rh��#��������)k�%R1Z����=ydn�� �;�
,��p�DL�������V>�;1��k�b��m��������YKm�4���oH����So�yD@���T!=��[�s�c�rg�H2Ruvۊ���!.?�����v1��h� �.sf�(n
�)b�0 �k,zz1(�3d�����[�B�X���"���M���n��]��0��|)��s*7�'(��bd_1���OkGEl^Οq���r�vE�v�E�U���JLq�\�Ŝ�zP?���17b��*�veH�!��g0K�"Q�cQ�?XlV�-�:Eܯ�_7����p�f&u��^�ڃ��J��`L��`'ZP�:� �DY�V���׮��[�9�&�[�`�����?���:��u�¼ ��o�
{"駡�<�2=�l��,E ��%X݅d��9)������������/����˷�=o��W�c��Z��8 >�����0 7S���+j#`���O����\�t3� .���_���XS�$Q�-����錨�GXRD���Ibct�'��)T󒴹"�L92�-1�Ǹ���4:��Vv��:
,r�0_Pi6�U���\d p������O& �2p�QS3(3H��g���#'�AM�,���&�;=��(��%oL)NH���k���@Q��0�S@�c|��
i�X�Z{�'���>�ڋ�(i�r���<�g���R��;��
��b�Hv=3��Os�~V��c��H9[k��[d�{�i���c[����*�Bf[����P~��-\���WY�
��x�mAz�f�s�$��=Ң�6�*�m�����5>�R�Z5�Z�=��!3G����EK�p�Z��
���b:�`���R>ƒ>�*�8��9O��d��xՁ�e�nG�D���R��w�et�����{�U"3پƪ�� ���X�x��ы�BB�e���4)sL^��@�+ޙ�tY��2�idG�Lr?'���	vQo0���Ӝ�x��|p�v�_�L5�:e-����	�`�v�AW�F�M��t���%0��䕙_I +�0*a�]���o�*؎���u�o�v�-ӏ@Kjr�*�,8��!A��୓ݓb��i1�"}t0���<��2	ˏ���8��2��KD
qF��x�����f#I��#7.��X�W|�ڿ*g��@X���avw��I
nw<���"��� d���i���f9�Y��<#с�]~��%?6�-Cl,eD K��@WɬD�&?�)./�w7[�-�6EC��)vلآ�<V�w�A��
58U,:ƗEN����c
A����J��|�n��5)A�u!��A�JQ�K1�~�e�ȸ�X����,?�yR{�mb�~{�J�6���#.0�Q�م�F)� �'?&�3yno�Q�X�ʞ8zx�Z�;���ݥ��>^[��\8.�x�� ڀ�C��/(^/���ȁ��~�M��X����Y��u49Qf�R���a��K
�A5J�m���j�Ŏ{>�Z-�h��<��7��� ��"�e�k�f����D��&�F���_�⌋��Q�[֥g�;�m �n˽U�h�E���'�=G����#B��誁�PT��"U2�䠄M�uة�5*)H��`�L%��B�2��@��:��Z�$F�@���[�CeJ�Ï��u�,�����'�M��
�!�"TK�7�jN�qB�fq���ϣB������x��|����X�����x2�7�dJ�����0v�H
I��KZ�����ep��;�!ePP�zL�m��q`/)jGϬ�fTm���`2rd0Ö��bx�e��E�2��l�]��-lxΤ���$e�(هzV�����`1���n�|�B8}�*�X�9��J�I���X�FD��O���nAgܤԱ���yY��F��mH�K��cA�\�ݥ�0eG��T�غ�
>hS:R�����ժ��#L7E���B��4�N^sf�A��a��?5r
Wм�͸�(��1�K�J�F�{/�8r�zM��T=�A��ӈ�.�^��,g�ߔ5i���WGM�j#�$�N�D=R��T#`I?a��x�ࣀ
[a[�{��==vұ�3ۺ��7��Ia?�LS.c��f)%&�M@>)�H�S�ŀ o��N[�(�0��c�z®�aj�<�����7��9�(��KF���ˈ��rk�A�����j�'{���4�Ѽ|F�WG\��^�N��Ֆ�@T�*띑���%(f`��~����6k��&�h�����ʰ2NF�]�FU��hF����	�	�;ϲ�Oڡ �)2~��:.��,� �r��@x&��ǚ6�fx�E$�1���EM,�����yl���Ɣ��`���s@����<W3����5��}E����b��ע�0�=�=-],K�15ũ��b{�M�{�%!=��/��בd�NW ��:ן�?�t�J��?�5`p���mb�E�	���Cn��$1�;}lJ�}*uc�eO\�s&���ҝ}�$;��F���:�����d�Ctqv_��{�?CHq����Q�s�e#<�ɔ� L�a ��䚡g�^ �#Q� ]�9���A��P�)ˑZڙ��a�M���}�/F�Y��?#3�k��њS�*gݽ1b�	�_��z_�as��"�j�Ζd�[�i��<�x�B���SF��	 KQE��M�WV�,S�p;o�G�kV�a�5
�yn�����z�aF�W�����v��%OTXP�O"5���M{���b�<Cp*�V�NY[��S��矯���� ��J�&���!���ɏB.=���e]A��^-)	�I�N��5$j���ݚ���B/��4��.��	P���v�}ؓ�U�@^N����m���
T�|ȣ�>:>	�r~$6 9���	6y�԰�Yyd�U!�֚8�v�����R���P�~���m�
q�x�?�5�	~����eTݾ��[�'���)>�4��f�n���\	7��D7����軄{_ tzP��X�`�0xA�av@��8)��,���5�O�w�����z�n�1n��T 6x���I�q����_@��O&:�3�Q��I{젧����{}���$����BZ�wHj~l��$#2G!U`d?6�0�F{?��
��Hi@A�"_���i��f%]��T߁��7@�7�(����H=ə��p�p�2i$��&����R+-E�u�(�r^��,�n��C_�d��ܾ�m��%��!�7�YR�ǃ5�+O�$n%�_�6m���f�2���6α��{��dŨ~�4(�V��B܏2����6f�XN�i���h�R��mf�-+顚���im��G�$����o���{b�ۺ�il��Ey��?`w(Ǩ���#w3�4�9B�.�f�`��O
���(�W�v�V�����/���<��|�ft��@��H�|#�\��`���E������F�-Zڻ�2�I��>��u����?��P�.Z��40 ��<��*/�`r�J����=�}ࠍ(����c&��
(�6��:�ɌU�/�_�+�P��@��7�;/�u��x_��=��ݟ8��z��ՍYNh3ݽ�V!�g�Q_������a�иËa�c����B��1fuk�K�i(6�˛�+��8Y�χ�R�2h���?$e<	���,��R�6�4"b��G��p�eJ�t�4�C|��kW�/��GbX�s���W��6����}@�ސᝉx�`��zU!Kf�0თ
�am_
X	�\��9��nv�u��wv��b���ح.l��s�;�O�
�D�y�˷����:�bш)��U�0#�HҢ�4.e��!>�կt���F*���r�^��w�L�N)b]]��i2c�Ɠ��O/�:�D�Y��Sf����0|)�ۂm�u�ʉ��d�B)I�;ժ"�vEk�*�,L݄��3�]�����HW���N7YF�9�৪� �k���MIB�`��P{"�7@X��w� @6gE{	Y�#0����W��x�x�-f��\����(v���a�_�in!���_9#M��m��M`�.��EWۂ��xy	G��,����#/K���0i]IR䛹����[y/j��nѭ���x� ���B�?%d������,TF�;oPZ��2�4Ɩ�Y�8H&yX]�TGu�Q6������2���YR�ؚ;��k�Q�������i��TV�WKz�VN)��9�}U�1�V�t56��j���J/�Dl�努��Ki�<�V��!��1�־��4e�Q�|�H�q�ԝ��382�}Z���i���(̵r9ʙ��$$��`�j"cI��UEL-�_d��c���l�P���lzK�}ݧI��v�ۣ�h��o�?PoJ�F��m�$�vu��$,=�Zn>��v�vBT���K�����Ay����iA2�{�]�}��?�?�DY��Tw�Xl�v>�6�F^*���>]��8���8;g�?��Ǘ�������-�����(t>�d���9�g2���2�J�S�-1�<Z���&��ү6���f՘L�G؝�oD�ɺ�*�]����ٮ��}���daA�E%�~�Z#��S#�.K�K�5��u��1�6ј6|�v����0`�R0W �B(�!�C�F��&^�7�gu��d�O�74�*c�~�=U:M������󌁜��( ��:.�u�n6H�	��@� ���^k�J4����sgw++�!z�q���1�\:�[�����M,>�&�~��̿�ó.A������D5d�y�=
�=Vrc�ѱ����m��T���M6H�0�W�r�siɌJ��)-��զ;����0x�,Ab��u�ꩽ�>�� �9��A�?�� ��V�M%�X��w�ᩦ�[�C�;�@Q�d>�s����>�f�g]��0m�Ʈ���
�� �
p��������; '?;��I.�i�BRN��J�J�"��١���A#�n��?��(�uD��\a�P>m_6|ƫF���-��z}<p������\c��b<��UO�IT��9Za����y��~*=��4~&��Y[k�˝+D�\O��+�R픦�W��dC
a�4�0o�/H�$3Y��Kx���|������،�����^�vt�6��zP��.�on����Ng���Y~�';�HF(J%�@#�پ�0|N�R��3�t��j@�ki�j��D�h�?�,l|�z�д�_��#���[u��Â(s��.�=���)�B�⁉n	5X�o�Eû,��`9>�~*���'לڰ3�S�����G~��erGKv�Ӡ,;9kl�M#5�>���'*B���"+�
.>{�JC�c��.�K�s��Sև��ȧ,���.Q?zѓ�Dd/W�uV�(t�]u<��X� �G.�N�e�4�BH%V �����7@��5�F�	��/q�L-��`�^�:�*��R�q��v%�"vW�><�J���	�y�g؆\���&� 
IT����C���X9]�22��Q�`�-��:���ҭ�~�S7 /��]Ww�3�x;��B�<y����|��"����f?��DV�^�L�Z� �'DG���&�)P+"��[������q4z�0�a�������^�z��%�����T�S�H�s޷a�F�;Ր���m>MV޲�O�ʫez����:�ɽ�_�v�u�a�/N`3sV�&}ט���| �E��-��e�AS�WK��7��B���5R��4�/�}'����Pk�h��@=x���O�#4��dz���:�*^�����wB���5�ɇP������_uK��������"��*�U�aǠo�A �L�!��E'J�%@��mDrQ��/$��:)y�HEYH�P`_��8U�;T��DaF�G#�5���0]#N�/���E���t�y<g�nX�'�I�oF
es�W��6��s,+ ��ɛp��}��Ȼ[HL���ӷ��oc�*@_��!"v�0�A����z�r�5I��砲�G�)�;�|�S��X_��G��~��G�@�)1��[P� ���B[���O}y3���L���h_�VI='4�A��[N���A����N�.�޻�*��6k�)B=�ܖ��N�n����u4����!Mk�n��|7/ W�t{�O=�)���>�����s+��m��H�.{��Z:�5��[iv�t�EI	íd>$�(���rO�I�L��4�"�C) �;�L9����B�S��\8��wi���2c���γ䐼�0��\�3ɑ�xW{��� �-��pA�#�n봏��nP�����q<Ӑ����0���a��s[o ������FO�7�J�׮Jvc-�{P1��s�Kp�i�	A���x�18*Қ!m�[���j�X&���7R�5�p����Ea�a��C��r��UB#�6Y���K��[�N�S}f����y7�ի������B���lGC��۝O.JZ\W'��¦u��ed0m���+��(���"�.�U�Y�myc͔���by�V�zS�����B��~ �/�
��Å�x��4U��y�b��`K�W�kh]�ŷ�؈�9�A�.�)+`O�Tl�M��uqҷ�������{q������0��?j���$l_"\8.�B�<�K��f������=�vwD.�����܋�M0i4��7��D\����^M��ί<Xh�}���@�X��=�h��ĳ�	�k���p�@�طW�+�OD3���|�M��w-8�7�^�WNOY_&��%��wY�>n{