XlxV64EB    fa00    1950ꗥ䞄;� !s�l:8���+_�\�x$�A��WF�on�l��Ź�
p]!�
���(�[?״��r��L��TnRI^�@_=Ҳ� ��9��J���Ҩ�b���	�O�L�7�=������;h�P���&��#���9!��Ju���\A��W3Ax"NT���!d�����0;�C�WS�^,Ł���T�t��ߜ�_f���='�x����OPMݯ��(��"c%�����	��h��=3ႆ�qyT�1���d^��'~�`�[�#��	U�&�=B��k��|@���Ԅ�;�mN�v_G��r�D�.o���}#��J�X�3��L�>}��Op��(�:�$��GS�"�i⚞�W
@�p��(��Z��(�f��y���'�����k� D1{$��0�>���	��h��EQ���P��>_	j��k]Fc�ƑE�x� ՞�h@ʃX�8z�pTJ�E����e����Brw����y�
�n���o{f<�B�p�Y�I��NYl��{�;*f]ۛu?�\ۙ>.S4�#�1v�(��Z�q�K)HK��(y��E�y��9sf���Ha�׵)�<t�\{�����6�o^��9��v/'���䈨/�6�e�o\T@Ay�����Ǩ�'���z��v�+����j	@�2���=,;�>
F��{;,�|Tfi�E�A�X��)������ش�B&Hɘ�a��
`ѳ�v���Eɦ��K�Lo��Y���!���.�Q��!�q�s��f::���MNA����אT^i�ݿ�g֤�0_�#�7NpG�(��݈�x�p�x*k��Q	zc�����%����jx�	�*�-��I����PHǒw����s��V�%X�/Ɠ0�@&ya��=�鐗	tk`F
��\z��G���ƪ�@(�4~��^;�Wp�=7��x�h��dXm�k��џ�f���bI/���xl� >��󂑒����b����pB�o�U�b_"16I��L/��¼�<?�\`鿢���8F��������#�&��4��¿"��[���!�Ldr��;⦏�k���e�8�fI?��/���V��(�\��dR��h&NO�&�SB�mV0���p�x��`��2�2�e��b������i���6?��c�j/�󙃄Y��	��pb�9�����U��@��e�QP��%�,2[V��iMe�8�m��/=­
����6l� �y3閂���1�r~�ٽ�������X��Ý��x[7���f�.�.�
�_c�c�lAS��l�[�b��Hܜ�,{jx]���g�2
���R�~D�+�	r���뢊b�eM6�h�>!Y	�\�u�Ů+.ך���H���O~(�:F�<FX��#�_S�6E|��|x:�%��������؟R�wV�e�W�i.��	��)n˔t��9m��</�8O�z���zD��B�����ܮ@�e��J��"��ܫ�y�`���I�$	]Hq��N�uG)���q"n��e��F\����#uj��FI��;�&��
E�s�t���O� .���T���e`���U�>r��������SMIضqu�/6���
'}4���	�]3��9����V���A=1�G�q'Z`�0ݹ����C�Ʈɂ�0�:x��Z��}l.����0��r�0Mq�[�v8i,`#��%W����x�����a��O�>(�T�����^D<Lf�;Ҋ⮡�K����n�R��(1`l`�a��g5�� ���F*����N��Be�� a�ܣ�����2��I��髏�ni�"]ݘ8�m����kMG���9y���X{�e@���,�M� x2����3�O��[��O�
 �cA�Up�m��-��#�h$�J������vɶ�D�V,�t�ׅyU�y^�Dr_�YG������~OgHNf2F�K�����`�eƞ����e��j�aK��80l�ґ�gHADg�ԅ�Z�����=��,	+@W@S�?1=���a�P'���d���ƂX��:� w���@��t��Gͪ+ٛ,eނf� #dm~δŲ��l�_>"���F0@� �����E�o{���.fm�(f��z�2�Y$�(q�Q���͹Ol�����K4�<��G�0k��B�݃T��+��0��S�x�K�w�P������>��i�:O�.���C	B�4k�R�8y\�b*4��SRV%��q�Oos�]���]�4������`z��axW�(�|�Ri������d���5=�"UOhil5E!�dQ��/LF��md��}C��"�O ��
�H/�Hg�e|����V����p%�w�c�W�|��8�ሶFp�Q�o�m%����4C���0��`�=��H[,lvV+>2c'�bLՃ���?<BUE��k�з2a-R
Zhx�Z�@N��~�/��n>�9m]����4�!�c�s稃�X�!�������* yz��i	�G�ٙ�9`��#V���E-t c��(}�q�R�&4:᩼�5qptcl�=?Q�����s��醀Η����An��@�*�5p(�y�}����HׅY���𖹅�R�ْ��T�_}��Ko.�_##��I��*#*���AXm��:��^���]מ��h���_��d4�7�u��H�n�5r�0��-h'Ԧ/�$�j@X��2���<0n��n���G��F���a�~m�ݶGH*��5�!��Uh�?���Od);����u��/�' !V6I'}��n�#e���v'�|,e�l`�D@�?X�G�?O�ǔ����4[��-y�wce�_��
�ǚ-��{Bȇ�5 �bpW��ݢ�M̪����&�~?(/a�Ł�v���k1)߆P�LZ��?�E��a,��Kl:���F�H�QSH�s�����ζQt^��,�!���zJG  �]�:�����X�K��lj�����<�Z,5������o�Kn��"��F�'#�R�\�3/�%��f�7[�̒93o6�"Y*;&g`Uݐ�"�dv�=C=/X^d8�[��v�A��f$/ij�Hvt[X��+�˳\2��s���1,�1�4f�ƅTZI�-l�y'O�(Ol,��8 �4t&S㏌���x}���G��k��D/�u�{��^��琸���q$+��z�u�߳�HG.	��ۛ���0ӕ��;�,;�!Z�l�)���"���nx�k�V1���� �`	=� ��3u�-(���Yx�+�D����[�vC�p�}iZ��W��چ�ͨ恎��=��Z%����Գ�c���oCm�P�S?!@*�M<��*�G�+E�>��&�(�ço��w`S)/+}�)�P,A=^�]/�]���Yg`E.��_r�lSRX���	�>���3$~ezV�0�BZ �7Ω�1��U�����TMw�Ķ�S���)��ݼ��׏gt�$��*`�ǿF?jV���<%`�p��i���A��+�w�'<��K��v��Y����ivP\�Kz�韲4+w�w��0��`}Q��ۚ��ڰ�<\N�R�;g1�D�ڋ�Ry�9?�����KC�ü�s�V�ۭ`��`ZIZ��f���PS=���g5�e��z�IC��Y׽�acj��]V��!��تCA#�Y�Z�3�I3Y��䣉ICD8q��I���w��G�Ց�w��үX��7���C	A��$Dy��Y�u����Np�0�\�����L�D��
��#L��݃�~���\�9��˯��)�`���ϗ]׀j��̣�D�2t���	��$�j���3��B�X+`�Z�SɫR�i�A���Y���6�����"��D��Zm�6�(OU��e���'���aWWY+*�<�wb�Y�fS�S�m�A5�����9� buB4��z|�辈%���^�bݫ��}��!Xd�� �}�5��jɱ`-���A�5��d������!y�%�w�h��n���f�x�a���5���4g�p^u�� ��F���n��@�V�-N������4�ٚ0�?d��B�c���
#�J����X�mt��Y�R'X����eM����]��(�'����r��ʳ�8׬�hy&z��dNޒ'�p�ƙcL��u��{�ȵ~5����T����|���$K7������{F��UTo<Nl�����Ըycbٹ�ocC�^�wh�B�F�N�����y�[!����r7c�0�٬���|dCX�����{n`Ҟ�C��G&�w54.Ѐ�HБ3��dT���H��~�,��+h4HjqQ�nr#�Dg�}�i ٪����O�Ёd�*H��!��l��	�������!�����{�f8y*4� j���Ǵ�u(����n\BC�RO��ʑ����b_�{Ąl����2�9�>�d����G���e���eZ��q�����F��b��� �+��&>��l�p04��z�$y��AhBA2D�d޽���*��nhc	�8㴂�r�C���׏w� 'C��|���j	ix|A���L��Ï�0�V��v�	bV"���B���� O�y�5�q"�8aTZlH_Q�X�5��]��R^��t��������	z� ކ$�������0����
ʲ
@�6�u�� �XĖ�59F��MZF��W�8g����TdZ�"���.P�!b�����*	���͂����~&Y�.NU67�+����9ƿ7�M# �p<
- �TpXW1Ee�1��`!Z=�V'Y�b�m;@=:QW����Fˡ6���*���L�h~�@O��Sʑ�nL2ċ�_��=�1$f9"�{�`p�$�FX@��M ���j܇���b�۩G�+d�mEƢ�U���^���8��tg��[�!s.�Gg OZ-�/|"Ԥ�,��L:!�J\�s^AX��/�&�pn[P�{�P���%8oX�f���'v�޷���zΑ�B���.�a<��_���sřĵC�-�x����?��O������`��J�o܊�¾Ʋ��������gą@�3��6�vuEW�B�a�ъʠ��Ec��}���J�&�OM�F:����/+���/�,6�SZCx�����!	Q$��}��R¸�J?C@��6,F��u�u���A�m������S���͊>��w���M���T/��M	���D��,�P�e9�+emKEl�<y�MX7�Ki�)�`|z��=r��'��	��c+�5��D�a���=
&�;,��Í@��ֱ��h�1�ұ~Ka��<B�ө
�$,�������qa�b����H�$�����E��o�a�l��7�\)o	xs%��[��jTT�x������]��D��YQD��p'�0 Yh,��ѻb���0]�9�t�!��(��̎y½�:1��J� v��K�n�'���g�/��:�1���������	~c�YC��ͪ�d�JkAZ'$��KXte?��ay�M��5�5�/���!��j'��9]��B�&���Nu��#`n?��}o��umQJ�>�h�G'��t��K�ѱ�6{�́r;�/��Tw��˦􃗨{�����~�A%B��J~lvlx�;���A� 2����-%5."�p�'@<����ĺ�(�[���xs�v��8޽�v�3�oX$�.ط˱s!)��5cl��q_�z+�r�. 
���w�m�<�$0w��d���FD�M�c	�@K3�L��P��g���$E��m����@��٦����3<����&�[��|�ki���T��\mZ-�~W\�_2!�{����*D�_[M /�������\fy8/���%J7��v~7VW"�!�ϒ�Q{_׬m���Ġ�M�Bam�sG%��l���la��~7Q�nc�e:����EV�4�[aUZԜ�P?Ғ�'=��&X �^�x�ZH��Rϼ��Q���DI|�%����H�s>-Z�Ha�%|��ގpH�u޾�0�Ɍŧ��!S���\��	��~��0���o�ޠ��j}�-{�pi�PS�ɕ�54�P��ԁ#�b4gv���A�s7HE�vt�/���W+�*A��۵)'��h�\�v[*��MH��s׭�l����fÑQi�;~��y"���;��҆��`��^�v1=|��F������7������?�3�Y�����u�����M��d�$ԫ��v?!��XF�F�!����x�5�lǈrX/Y�Kx ]��|B\��DnS"ޒF֗(��Aą����J�u! ���I���6q�yX��5�ɥ����u�pۤ~H�Ỡ�����H� ���N�H�S��3nR������X)t�i�0bm�6�`Wi�{�۷T�KإG�"�8ӳcq��G�	QN9u;K�h𛆤�X�XlxV64EB    fa00     700ʻlra�c�ʈtPx����N�DI~�����>S��,k��UpR�T̎�@-�o1�XЉ )�n̶�(`&��Y,?�Z!T�\���?��|�MҸ��.�6�
$�TY��������z?z��^��a0�X�S|-�NZ�J�R��7ՠ���V�V��Kp�a��]3i��f�g��$0��S�H��o[B�gt[[��	���mb��}��a�gж\��4]�Z&�Iᇾ�x��?�){'��]�yL~H�x֙Lz"�&���4�"Kq͗�'r�ĊF�yE1��3��@��j��J~���~`�謲L���:=�����p��nz%��$�?�K&��i�pA��|���NPo	�.�G���H���te$��c5^-�E������7\�mDS'�yl�y��8~���˫$x�2�$g�a6�۸�$���@޶ҏ�f1X3Ǭ�:)ʤ�|���T4�D;Q*�1
{X@����܁	I�u��"t,�CЊ�gS+��1#K�PR�B�~ۻq��}�8���{�&P�W qʨ_�/,b�}�Lif�u2�FXIa]�3KT�v�>~;o�v1m!O�$'�y8��+k+|����e~*]|��)�)@�Y��4�����b�&���JU{���#�͇��H�����ሺn�D�yq,�>������,R	J��>�5�ߣ�?;��u������v�7E����+o?�'����8 �� �^���U܎���O��g��!�+ך���=R=%��G����1sy��f�V(|(�H7Q�wA����طt�K&��,�W�I��m�_�}�(�>��?dr�������$�Wv��s��.y����kԸY��e-�2���t(�����mhn�S�IlAծ?탿��B��u���w=��=�E�(b(Љ��o���f(�"���K�M�
0��&eՒd�0g��[Oz�'�.Ǔ� a���6��*\(�0�����rG[^M�SE`P0��6=yk�0����V�j0#�<7���k��(�s��׫��=D����0��R!�Ijd�r#��>��w"(����/Q!h�!�'�Z��k���"�mW�1�r�u�G�+(\H�u����A]�s(`�'�;����۸bc�z5�?�ø07h�G��/����I�z1���e��[v�!K��fN���	6�u�,�  =5��Ԑ���4���؎M��b6�Mȡ��[1?e@w��ȋL�� m��=O�ůxyB(��<��*��⌇M�q{׺͠����2��S\���YgC���3��՘˼Gg:rO���{>��:3�z�p���g�t�jb��|Q����љL����e�CEGH�����MQ��P%�S�G�8�<�qɅ�l����.yq}��<,�N����V��=|���k�ND{ب�/��Ra���u'�6�2Kl�H�]�y�f����P�)B�ło�x��Y�������3s���R��{��-�4���m�.^����FO��8��������Z�Ep��#wf+��B�m0WɝrMg�e41�4��5���ђ���<�����QU���;H�B�wܴ�u)��m�����J��C�#g,gv�>�D�$��w</&hD�o�}]1Q��+�t^����
̇F��D\�v�7ԟ@؞Q��P?�zJ1��|��\�S���چ�Q&YÞ).0�'�E�n;�gFX�/:xmb���o����Ļr�/!*~Ek�Ё��v�S�\�*�m�����XlxV64EB    7d01     bc0�c�a�o.��_�B�)I`ι��2~sGm��������F��K��wI�&�1Q�����O�	|�5�t��wYKL�u@a�wo��>��hF��8��u���l�%
��Eޅ���h�l��>�zoB��D�~W@U�޴Q�I9>�Z�e���DH�$"�+�j6q���u�g�h����v���׿���*�VN��o'��=�~��y�&
v$0��5��l'	z|�a���L�Ne�@7<��S��6��G����5&�7��1���:���Y\��S�6�?��6���+�.�(Q��b����uX��A�5;�;�u	��ܿH\b�0��9 I�n��!v*���E9R`�����5o���{*du���ArW�D��J�F����<d��긹4I�A�_�$6�9����5�b�!@���2'�k �c6VJ�Һ�N���8>�	E��~��h�B���s��ק.�B[Q�ݡ��H>��:�q�=1���2�H���,�յJ����[/����-?��t�ܾ�V5{�^���=o�q]t��dJ�#�6M63�f��+j�Ad�&\di3�����?D�^�oB�����O��n��}��T��B�9k���!��tDN��ב�'E�p���@1L������y�w�v!���D�lXg�����B#��^x��_����$zf݉|:�؈<�E�a0V���Q��#὏�p�j��L$:�(i�����|���@�y&{�C�zA�
����Q��I�_٧�ڡP\O؈]`C��S��߽�NȪˢ�焂߶�a��wy =�0l�e�͓jưG%eA�$�D��hlWK��̢q٭G�:��{������yȹhe:e���T��z��#��F���V)�s���:���*���)"��������X�!X���wq����>Epp�8� 7�$c9�+!<n�O�)C�7�[fk��0�,����.4���q4�~�����"Ts!X(�2��	;&q1z�`�WI��VN�2t��+�G�Z��JԵpQ�H5P��j7��]��ZR���SB84J��hq�+�&H���#�H�#�j+}d˴;;�nLn酷���;��OTC�����C��N�cV-"�[�
����4ci�D�a=g��=�s�2C�kg��\�q�j��j��w,>�%���Un����_�P��VC>&rf�JR	�p?,�E��7����c5;Q�z�&	c�b!5f��(~��8�Ґ��1Orf9��q	�y�)�f�Q���D��	`f>z3�r�Y/�x�剥f�b	�yA��}'��u,|NBiܐ��8�<�8�-c�AЀV�ե/��tT�\&�ξƔi,K|<��MI�[º>ý�)E`�l$�ۼ{C�+�P�6���!��u'�f�<�6˘>�$����nώd����aҭ�:>��Fu�[�[����҄C55���<�"��Bxmޕ���I>�B�2��鎤";���a�+'���Ѿ�s�)�dw٭�.pm��	ߙ�\����Q�Ϲ:6xl
a��<���Nۣ��NϷ7U��̭���Z|;�zM��F��Wa��Z�ᜄT��ne:��9�L�_��(_���A�N�͊�p��zG�A�g�b�'�3gh�21��y /�L!�ē�����v��� ���I���X>=����h��S���mdk�=l�����u1,3$=
��P�Q~��/w�;��,/J��.���V52��]���������u��FˀjĤE+s���t���~� �������c��s.=�\��T�'�7G#�q�<��f��ݧ)r�-�A�P^�*^qn��1LOu���)���[��Ƶ 쩰}!��L��=/KV2AƖ?�'(WO �����w�歫L�{�����3�A�ϧF`�O��9u$�}��jc��y��^��:*�8��W�\�=�[���c���N�U2+M�����cӖ� ���x/���a�����_>����I2q;�E".L���g���<Z|m��qS��)`��_)�j�?�ź�H�C��X�f~}�	nɳg/y��;��MD�d����X���/ߣ<�1sWO:V(Pi�3�%�Vc2+�&þ���r�GUC����>?���r�[�v�:��U�H#)���m{��� >5"���Ə�Rk��>AgF��^���֘6W�;���񁤣_�⸇ⶎAgz�8���b�k�ϪFa���{�i"#���g�'��Sa7t�5d�L��}�̈́4�o6�i`Im�Gd��e��*:���ʧt7�5�b�V,7g
��C�ݍ�j7�:��Ϳ�z�)��:dE�Ŝ����k�<�IG�.2�c��2t����D�"�9���U��H'�D�E���:��lK\���)�!�ap�'�����0|ђ�"����������_��i��.��;���}ѭ����Z�k�t����{I���,ՠC]�Wu ]����w�V�M//��׭�ď�I��h� �k�Kr;�@��݌�%����^���.&Lv�"7?Y
�ee�/�5�Y�&�Z�L��`����P���bφQ�%�k�dS\��	(�`���\bmI$��*�՚��6�s#5�%.���W�I��k-c;��th�؈�hRP�I�o�i�8����DZ�w's�^��d&lc�����}=���:�8Y�g�kNc�ݯ��N�p8��5��,��0j�2y(�"�4��F!i50�~0TQ߷��d�Q==S�9�?� ��1��߂��������O�D%��n����qsA��3E�~0cOQ]7�2چ�[λT��p9�i�녕�n5P�ƅm��e�r�ΦN��h�T��QئcD���K�v�-��ʗH��&B�oD�t���(<�_!�1����J��H�B+��RøлE*x�w~Δv��Ppю(��R����-ݿ����*~G���6