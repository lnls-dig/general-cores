XlxV64EB    6dbd    1650U䫍�ޝ�K?��_�(>E���U^%Ʌ���W����ԍ2�jSg��偀8Y��>�{�5�������<'��Ĭ�*�G�!t�����n�(&�SޤdV`F3� t�{Q@��,�Ү	Ep����@����mшhH�6��&QE�Fi�@S�F7�Z5�0>A�i����3�R%�R-a��H��(����>.�~��'$[������q��vDl?��_dѯ�	FT��)�e��y���fz��k��߈�ǵ�a7��&�[�.��c�3S�P�G��n<$�7a��x$<�.��W�����:>��YT�[�O^�xP�ݟ�;�vI��v��V�!��iOcY�����h8�1u���[�'�҉��R0�Ř�4򟩏�x"~�de���4�}�T�]�p��S�(�Ճ�=�l(�2�8FV�Q�p�Ԗ%=5��-�����5��Kաx�g����;X�yF�ao@V��wĀx�
����sV"�3�� ����$��|�����1
l��I����t�>��	nJ��$*tXg2C[���r-���X��� g��s]���>�?������V�o��-���k�P+�׫{:$�%�񓥉�S ^��<�(�|g�u]�^C�����ߠ������w��̹����Ƈ��?J����J�������F�\_	�	���,�ݶ�}&�YbA����\�:�V����׌L�?���H9b����]V|r;S�����7]���9}�9��KO���8���8�;� P��^��0�D�kΗ���g Qy����1W6q�o�f��L����SJ����u�;(@v��c5?����P���)���|�XWu�ߪޱd�b�џ����?�����_��Ȼ��f뛩���+��`���+^G)�����"�����g�c枮�y��&��F!�$��Ⱦ�ޣh��6��S���_\}��D��b��h8a��%�W��ĺ̏D|���؋ ��8!f㫚-P؃�s=�� �0�U�#Y�>��A6�%��h "��j�6z��v�w�B��愺���M��+��ԤkVAx���T��y��Q/�t�z4���	n�p�1� {rϊ���*�a/��&t�5�����ߪ������b��`�`������}���v�ETW�;}�ҿ��]��ыmV�y�s��BT��OXr�� t(A@W,�������� ��"G D+{����/.v�Jv������Y	(�v��ZL]頢\7��;�^6~�����
���b��[gg�ե�>�g��c"mޙhL#q�Gy��Zz �����z�d�4�aD�,�D.�R�:5ͩA�ßĂ8pd�y�$XO/<?�P�?�V��CLF�B��Ӡ麔��84�QC�{�+ +j_� �X^�ۢR��a_�
��L�p�4�2x^<繲�};�󤘬g�M�"�o�:���}vEY�V>z��,yc��I�F�q�+��*&��%��)	� &u���R�,o��� 38#���Jyۗwހ����'���l�T��J�����)�h�ݽ5��N�4��kT�D��VΔ�n�Z�䴏��>�pf���g�$f�?�:�,@ �.�����Q�p���@ *�ցώk~�:��.=���kb_�h�ͅM�`X7�����!��g� :C�Z
28vDMyל�1��&�6�c�wDHQ�ˉ�'�F7�DL��};N�|.Pm�]rS��6�����L�s��f;���u,�>��o�k��	.�n.�O9m��s�<Q[)���~�n���}g��c2�".�}�)�q�o�?�$��A	�|�q�05�M���/M�Q���ܩ6��ru�˦Q���K�V*@س��!Y
!��~;H�*/Sx���^�F��O��e۠��zl�L����$�Munڠp6�)[Yy�ݠb^�Z�����*dЖ�$�H�_ę� 6 ���Qzl��\ �WY�r��qx�r��e�_��\z32"��;r�O�Kvn����_��8�;�` ��t������z��kH�C�$�_j����#?)+�S�A�R���������^5�l���R)��ҕ7�G;6�HGLf7u!}���V����+��#�U�Ә��AӞ�6b�j��&��c���Pg��Հv�{itU��ρ��?�lL��T\��uXR}���#V�ăb�<��˞j�B�=~�f���2pG��|��4,�V�%_��<��p�VV�"C�ٯ:��i�Co������25�?H<���p1���Fv�!	^I��H�w�$(���A^>����ܘ���8�Il�`a�T/< �C�r���?�m������B(s{/���JL�n_�$;���Bn��2j^.���Z�77��8BU��~�AVX+aa�-��v�q)���y����,1���'�ʇ� s��&JE@J��U�GP�2��e��B��W8�ޖ�6}|�h ���T�#�J��� \,1b�R�23%�&�����MD���x��R�y��-@�oT������h�7�w9B���M�S��C���f��}��^���t/i���:�����]澐k��H	<�z�v�E$6pE�+D3�[d]@�tE#0ER���b�/RgTu���:������M��_�l��r\=����uQ��.as<ps��~�[��X�+[f�ګXx-`��?�����b��3PH�����	�	uU�󀒆]6�5_
��u���ۋ���_�L/Jɿ-��KÀ^�1��,���k�&���Jf����B�(6k�C��������n|v���etAq�
�����̧Q�<�6�,H��f��T�0g��~��&��p�&����>-L3R=�Nd�����z�T�A�j*/���$r�/�L��&��<IhKu����[�@/����?�Ќ��3��-�����d�����o@lg�B���t|A%u�Ηq'=M$R�+��	�f}����KGO^ZR���@P�if�#ru���+37~�$�U�]�>��!r���jo��JٟP���Ҁ��J\殒 ���7^��Q�����ʀ��&fB`]J���cí�f���{��{��ED��&���Ƈƫ���E�x�1]��Wہ�,H��:�JefG� _ٚTϦ$�f����9�,��Y���ƴ�B^����XlZS�	��Q�?~$Z��I�R�Y8�¨�A,N�xm�|Ssa��lH���4��C�]�n(���C�>0�I+BC���t��4#6�2A
e�=',��KKƢ��+@�7c-)�c6G�\�8�#�6�ʸ|��V��R6&P��ݠ`� ���fF�F5�!� ����슄��T
"�h��4���[��QgցǶz�a��L��2�ɇ�9\+��Ġ��r�����b�y��]&u��b�*��r#�p�n�X���h��`Z�l�˴��r�U ���&<�"��蜅� ���
 
겊�<�0&�Ƭ��ϰcp-5���&Z�枮l���i���ì3�X�g_J��x)4�<]bc��nb&���`��'�3ʡ�a�?�D���p6�rgb����v7ǻA�0����Qՠ$��'�bP+=�˺"�&�L�8" � $GGL�L#��!cC �Wy`��*�v�hd2���E�3U��<3�w�y�D&<ɛ�t��EST+*=��	��ؘ&E�\�a	Ӆ���"�����r��v�i?>��,�i+�F�Z(Q>�m�!~?\�'j���e����P�n=�}��a81����2x�f�0���5�f� ꭤռ�h�cVQ��[�U$�
jBӒ�ܳ9ӲվL �W�������֎�`B�=05�:��(9�r*N��t�`5�D�_�ASn�|6ׄ~Gtޝ�_��L��Z �s$���F�6��O\�L{�Drm��B?f9�3׫��y��Jn��,�y�ՙ�]�keINB��I��P��>Vl�N@��7x~���GOq�T]�M��m�˯vӷ��Q"g�m����/��p��y�����*�F��-��Q5�Gӥ�P�{3n� �T�V�����y���V�7��`�ʀ
\b� m��Nђp�r��z��w�z- �v;���¨�\�i��az���Dh���$q|��kPLGZn5��,s�(��CzB�Lo���.�����*��=e*e�6E�3����R�
��O��:cаy� �S��*}�0ӊ>����{�3�y��3�@iuG`��`��{�E��V� �q:��ܱdƢ>;w�"��]�+<¿�2�j-�T���4آn�艹��fd�.^J�!y>,�֞��4��gtg��g���%0�fO��~s��A��m�꧞"�t}�Ҍ�m��x�� |br�jx:+|�l3�q��&
� >v�m��E�tĂ�mǩ����i���jp�V|8L,��DA�&Z���e�SiŖ�M[NԤ��{���^�X���s!>�T{�H˨�G�C��B�7K�0u���GG��r.�bn�f�e55��P�t��=g v-f:�pz#�ҤHOe���S�/N�Q�6���h�<�7A2Z�`�?����>��]B�NK�1��OF�Ss[��c0��(��YvrC����ڦ�cDSDT>���
��[�T��I�C c��R��Qe�̾!Ӎy!5k��@6�q?�MY/��,�/�h��}D�HH
�}_H�ҵͬ'ӭ|�������!�I���In��Z+��՝�L�+ipF��Lq܊��ܦ���]'Cf�������qQ(W�E}j��c#��)�V�2���h�,~��-��ف� \���'�c���A����rK3����w�kw����O���NXq�5i2�,(��у�@c��+���Шo��mm�	��F� �e�XL�(M�-��3ȰiS����s�"�ൃ�u���~T�g�Л˦�!��ynDRK�p��0�j��/8�B1/:pC./����"�gZ#{�i�`�ֳ5���N�|���!ɦn�P��ȵņ�E��y2�h�O��5������!�7^��2�9�j|���a8���}��-�P˜$�8��%X�Z��Z�:�� R�\�y��6�?B������`8R�2�c)Ծ��R���=i˞���v^I�v�,���e6��t����r�$�J1���2�K�*b��C�t&\yT��r�@.SI;�
=���ͧ w�:a����_�KO�K+>��B���D�xU�V]pC=�ȓ�Y��SLD�B����˵h�rf�ev�_F<Sq�} ����;_�u�}v���s5���|�dAc��8�´�b�R;3Z�1v��V�i2H���z���7�V�{��c��1ⷞޏ&M�3ۏY��(�%�>�E;��:]�@�1�G��8g���C{�#� �CH[��W���Y�r,��
J|t��x[('7L)A�؃I�D�(h�e3�� ��G,8+g�6��7�y���B ��]^��c��E��6�� �S�!�倀�w�f�$�1��|�Й�w>�0���D{X�[�!���|��ɭ�I{�Tma����"7��}>�򍾛#�t�~�"�������o��b�Z��s�3�P����pӈm���F��٤BnM�����͎��Z�0
긧