XlxV64EB    1b42     980�&�����;q�tP	Κ_��Ph,��lY�����3u'�ܳ��s���0��y��<����@q���G�����uC�;ж��3{$K�r�Ky&�����W�]q+`�Zs�+sw6^H)|e�;��,0<3dF�j����(C��pO`T��؈�^�c�[g�ϒ�9&��F��.�[J����x<jm�N�0#�,�3����~P����2�\��Y�5�z��ֆ���=�"/w��|���Ot�v����~t��̾�R�qc��,���22��!s+��C�w�X���|<��/U.U��dOn�H{�\c>{0��GA��C���Y���Y�x�f<���ǓXv����]���S��z����R����<����M��v��qVlSAX��+�z�s�KR$6��p�SZ��ƴa�j}�����y���Ѡ���	Ivc��z#=8�D�۶R�^x����`�*�U��Sv	������9���?ҵ ��O&��hs�=;�|�jgQ
b��+S�ơ���EjT{?����\�L��"q'�������U��^2,r�WC������fK_Yw�����iP������˟��:�a�)$[�b.�Xz��N�b����*��.��f��S�_�͑�'=��1qmW�����	��V`���j���nþ�^�]̀/�m���6<{�f���4�ƧOy�D}[h�]U�ۥjT�ţF�*G=Ŧ�p���0K+k|��sWrي{jr'z�`�-dv���P��(��|b�����/qFb۠����&����o���3H
0�c0�|.���������.�}�]�ҵ~"i�I�J�wnHk�cL#ȼ�o���o�53��IE�����t.(@8^�6��ٛ��E��YT�8#~�-�(�_S$���Nj� =Y�D}��|��D3ېo~`���v͘RR/�{�ۢ��v��<"�jy��-e4���αU�́�"��j�9�N`Ǫ�{�!|�6٩|�������ǃl����4�y�

�_8^�C�3{d����`��vX����=Yl48���y(��¢�vؓ���
��?�;ne�Vkɭ! �iA�n�nU��F�f$�MXF�+5D�Z���_�Gh)��J�M�dZ���ž#�Wc&������g��+_���#xC����CiV��v��.Pw@�Ǘ�����Ҧ|wB����c	2O�u>�e���D:�R�W_����U���'�F�H4�ӑ��s�@
6���`��S�SU��t.�nT3V=Lo����-���!]*��g�p#䯍!�BSU��p�	h �U��[ ���U����}h�ӎ'6��1b�C(�W�?%9�F�G	�_�;�Bb��n���Ixs�;Hh8��G�Pƞ�AN����{R���~�Z���
��d(ϨQ{���'?����z�4�"t1C4���C�Цu�<�M�z��I����E�6�8��Ƌɩ�t]����BK�|�Ȃ��ڗPQ3����偭[oc�M�|�Ś�^&�a1�^�L�`��
�{�b"�5$�p�{��~x�A2n������>.�í�p��{�hn"Moc��bӀ�������+�Ն�}���u�\]�V{�'�����C�`}v����噶�~�{*c��j�Y�.�QO~/p��Wd�K�D�GR�q�&�Z�i�s����T0�9�૟�V��򲉗�"�I�]\_�B��5`�Y�"��iW�O`��n��js�؋��_����~�D}��t=����L<LVu1i���"���!I�)�-kϭIr�x���?��Ta�K�t��K�/](;���P��Q��d�"+zG��^k�������?2�J/����,�l�XW��,�.Vo-�R��
���ͧ�0|�IP��Y	՗:�?� ����p�)��>����d&��3��2�/�o6�ػ5m]_b�ۯ�p��P���G��],¡�����T!���B�� ]�f�8�/�T�e�������E��WۅE�'X~���g� �qB�e��C���Q$��/�j6p�E8 �0�5ժ�����/��^�l�&��<(�RW���K��M��/�-@H� 9ٰ���fš|3���-a�;�S������BF��q�"���SNz�0L��w���AF I�B�A6�js��{����P�[��s����-����é�d�y��N]�B2��g[f%��Oh�in����oG��'��_�&l*>�Q(����._�@U�t��e��J8}�k�x�ƃ���c�D��?�lH.�f.;66�;��@ޡ1:٦���R�H˒�Mؙk��$`a��CQ~.�#�xe��s�h��)w/�Să��Mc���)���a?�&f)�H�,��dˊ0_���u