`define ADDR_XLDR_CSR                  4'h0
`define XLDR_CSR_START_OFFSET 0
`define XLDR_CSR_START 32'h00000001
`define XLDR_CSR_DONE_OFFSET 1
`define XLDR_CSR_DONE 32'h00000002
`define XLDR_CSR_ERROR_OFFSET 2
`define XLDR_CSR_ERROR 32'h00000004
`define XLDR_CSR_BUSY_OFFSET 3
`define XLDR_CSR_BUSY 32'h00000008
`define XLDR_CSR_MSBF_OFFSET 4
`define XLDR_CSR_MSBF 32'h00000010
`define XLDR_CSR_SWRST_OFFSET 5
`define XLDR_CSR_SWRST 32'h00000020
`define XLDR_CSR_CLKDIV_OFFSET 8
`define XLDR_CSR_CLKDIV 32'h00003f00
`define ADDR_XLDR_FIFO_R0              4'h4
`define XLDR_FIFO_R0_XSIZE_OFFSET 0
`define XLDR_FIFO_R0_XSIZE 32'h00000003
`define XLDR_FIFO_R0_XLAST_OFFSET 2
`define XLDR_FIFO_R0_XLAST 32'h00000004
`define ADDR_XLDR_FIFO_R1              4'h8
`define XLDR_FIFO_R1_XDATA_OFFSET 0
`define XLDR_FIFO_R1_XDATA 32'hffffffff
`define ADDR_XLDR_FIFO_CSR             4'hc
`define XLDR_FIFO_CSR_FULL_OFFSET 16
`define XLDR_FIFO_CSR_FULL 32'h00010000
`define XLDR_FIFO_CSR_EMPTY_OFFSET 17
`define XLDR_FIFO_CSR_EMPTY 32'h00020000
`define XLDR_FIFO_CSR_USEDW_OFFSET 0
`define XLDR_FIFO_CSR_USEDW 32'h000000ff
