`define ADDR_FPG_CSR                   6'h0
`define FPG_CSR_TRIG0_OFFSET 0
`define FPG_CSR_TRIG0 32'h00000001
`define FPG_CSR_TRIG1_OFFSET 1
`define FPG_CSR_TRIG1 32'h00000002
`define FPG_CSR_TRIG2_OFFSET 2
`define FPG_CSR_TRIG2 32'h00000004
`define FPG_CSR_TRIG3_OFFSET 3
`define FPG_CSR_TRIG3 32'h00000008
`define FPG_CSR_TRIG4_OFFSET 4
`define FPG_CSR_TRIG4 32'h00000010
`define FPG_CSR_TRIG5_OFFSET 5
`define FPG_CSR_TRIG5 32'h00000020
`define FPG_CSR_TRIG6_OFFSET 6
`define FPG_CSR_TRIG6 32'h00000040
`define FPG_CSR_TRIG7_OFFSET 7
`define FPG_CSR_TRIG7 32'h00000080
`define FPG_CSR_FORCE0_OFFSET 8
`define FPG_CSR_FORCE0 32'h00000100
`define FPG_CSR_FORCE1_OFFSET 9
`define FPG_CSR_FORCE1 32'h00000200
`define FPG_CSR_FORCE2_OFFSET 10
`define FPG_CSR_FORCE2 32'h00000400
`define FPG_CSR_FORCE3_OFFSET 11
`define FPG_CSR_FORCE3 32'h00000800
`define FPG_CSR_FORCE4_OFFSET 12
`define FPG_CSR_FORCE4 32'h00001000
`define FPG_CSR_FORCE5_OFFSET 13
`define FPG_CSR_FORCE5 32'h00002000
`define FPG_CSR_READY_OFFSET 14
`define FPG_CSR_READY 32'h000fc000
`define FPG_CSR_PLL_RST_OFFSET 20
`define FPG_CSR_PLL_RST 32'h00100000
`define FPG_CSR_SERDES_RST_OFFSET 21
`define FPG_CSR_SERDES_RST 32'h00200000
`define FPG_CSR_PLL_LOCKED_OFFSET 22
`define FPG_CSR_PLL_LOCKED 32'h00400000
`define ADDR_FPG_OCR0                  6'h4
`define FPG_OCR0_PPS_OFFS_OFFSET 0
`define FPG_OCR0_PPS_OFFS 32'h0000000f
`define FPG_OCR0_FINE_OFFSET 4
`define FPG_OCR0_FINE 32'h00001ff0
`define FPG_OCR0_POL_OFFSET 13
`define FPG_OCR0_POL 32'h00002000
`define FPG_OCR0_MASK_OFFSET 14
`define FPG_OCR0_MASK 32'h003fc000
`define FPG_OCR0_CONT_OFFSET 22
`define FPG_OCR0_CONT 32'h00400000
`define FPG_OCR0_TRIG_SEL_OFFSET 23
`define FPG_OCR0_TRIG_SEL 32'h00800000
`define ADDR_FPG_OCR1                  6'h8
`define FPG_OCR1_PPS_OFFS_OFFSET 0
`define FPG_OCR1_PPS_OFFS 32'h0000000f
`define FPG_OCR1_FINE_OFFSET 4
`define FPG_OCR1_FINE 32'h00001ff0
`define FPG_OCR1_POL_OFFSET 13
`define FPG_OCR1_POL 32'h00002000
`define FPG_OCR1_MASK_OFFSET 14
`define FPG_OCR1_MASK 32'h003fc000
`define FPG_OCR1_CONT_OFFSET 22
`define FPG_OCR1_CONT 32'h00400000
`define FPG_OCR1_TRIG_SEL_OFFSET 23
`define FPG_OCR1_TRIG_SEL 32'h00800000
`define ADDR_FPG_OCR2                  6'hc
`define FPG_OCR2_PPS_OFFS_OFFSET 0
`define FPG_OCR2_PPS_OFFS 32'h0000000f
`define FPG_OCR2_FINE_OFFSET 4
`define FPG_OCR2_FINE 32'h00001ff0
`define FPG_OCR2_POL_OFFSET 13
`define FPG_OCR2_POL 32'h00002000
`define FPG_OCR2_MASK_OFFSET 14
`define FPG_OCR2_MASK 32'h003fc000
`define FPG_OCR2_CONT_OFFSET 22
`define FPG_OCR2_CONT 32'h00400000
`define FPG_OCR2_TRIG_SEL_OFFSET 23
`define FPG_OCR2_TRIG_SEL 32'h00800000
`define ADDR_FPG_OCR3                  6'h10
`define FPG_OCR3_PPS_OFFS_OFFSET 0
`define FPG_OCR3_PPS_OFFS 32'h0000000f
`define FPG_OCR3_FINE_OFFSET 4
`define FPG_OCR3_FINE 32'h00001ff0
`define FPG_OCR3_POL_OFFSET 13
`define FPG_OCR3_POL 32'h00002000
`define FPG_OCR3_MASK_OFFSET 14
`define FPG_OCR3_MASK 32'h003fc000
`define FPG_OCR3_CONT_OFFSET 22
`define FPG_OCR3_CONT 32'h00400000
`define FPG_OCR3_TRIG_SEL_OFFSET 23
`define FPG_OCR3_TRIG_SEL 32'h00800000
`define ADDR_FPG_OCR4                  6'h14
`define FPG_OCR4_PPS_OFFS_OFFSET 0
`define FPG_OCR4_PPS_OFFS 32'h0000000f
`define FPG_OCR4_FINE_OFFSET 4
`define FPG_OCR4_FINE 32'h00001ff0
`define FPG_OCR4_POL_OFFSET 13
`define FPG_OCR4_POL 32'h00002000
`define FPG_OCR4_MASK_OFFSET 14
`define FPG_OCR4_MASK 32'h003fc000
`define FPG_OCR4_CONT_OFFSET 22
`define FPG_OCR4_CONT 32'h00400000
`define FPG_OCR4_TRIG_SEL_OFFSET 23
`define FPG_OCR4_TRIG_SEL 32'h00800000
`define ADDR_FPG_OCR5                  6'h18
`define FPG_OCR5_PPS_OFFS_OFFSET 0
`define FPG_OCR5_PPS_OFFS 32'h0000000f
`define FPG_OCR5_FINE_OFFSET 4
`define FPG_OCR5_FINE 32'h00001ff0
`define FPG_OCR5_POL_OFFSET 13
`define FPG_OCR5_POL 32'h00002000
`define FPG_OCR5_MASK_OFFSET 14
`define FPG_OCR5_MASK 32'h003fc000
`define FPG_OCR5_CONT_OFFSET 22
`define FPG_OCR5_CONT 32'h00400000
`define FPG_OCR5_TRIG_SEL_OFFSET 23
`define FPG_OCR5_TRIG_SEL 32'h00800000
`define ADDR_FPG_OCR6                  6'h1c
`define FPG_OCR6_PPS_OFFS_OFFSET 0
`define FPG_OCR6_PPS_OFFS 32'h0000000f
`define FPG_OCR6_FINE_OFFSET 4
`define FPG_OCR6_FINE 32'h00001ff0
`define FPG_OCR6_POL_OFFSET 13
`define FPG_OCR6_POL 32'h00002000
`define FPG_OCR6_MASK_OFFSET 14
`define FPG_OCR6_MASK 32'h003fc000
`define FPG_OCR6_CONT_OFFSET 22
`define FPG_OCR6_CONT 32'h00400000
`define FPG_OCR6_TRIG_SEL_OFFSET 23
`define FPG_OCR6_TRIG_SEL 32'h00800000
`define ADDR_FPG_OCR7                  6'h20
`define FPG_OCR7_PPS_OFFS_OFFSET 0
`define FPG_OCR7_PPS_OFFS 32'h0000000f
`define FPG_OCR7_FINE_OFFSET 4
`define FPG_OCR7_FINE 32'h00001ff0
`define FPG_OCR7_POL_OFFSET 13
`define FPG_OCR7_POL 32'h00002000
`define FPG_OCR7_MASK_OFFSET 14
`define FPG_OCR7_MASK 32'h003fc000
`define FPG_OCR7_CONT_OFFSET 22
`define FPG_OCR7_CONT 32'h00400000
`define FPG_OCR7_TRIG_SEL_OFFSET 23
`define FPG_OCR7_TRIG_SEL 32'h00800000
`define ADDR_FPG_ODELAY_CALIB          6'h24
`define FPG_ODELAY_CALIB_RST_IDELAYCTRL_OFFSET 0
`define FPG_ODELAY_CALIB_RST_IDELAYCTRL 32'h00000001
`define FPG_ODELAY_CALIB_RST_ODELAY_OFFSET 1
`define FPG_ODELAY_CALIB_RST_ODELAY 32'h00000002
`define FPG_ODELAY_CALIB_RST_OSERDES_OFFSET 2
`define FPG_ODELAY_CALIB_RST_OSERDES 32'h00000004
`define FPG_ODELAY_CALIB_RDY_OFFSET 3
`define FPG_ODELAY_CALIB_RDY 32'h00000008
`define FPG_ODELAY_CALIB_VALUE_OFFSET 4
`define FPG_ODELAY_CALIB_VALUE 32'h00001ff0
`define FPG_ODELAY_CALIB_VALUE_UPDATE_OFFSET 13
`define FPG_ODELAY_CALIB_VALUE_UPDATE 32'h00002000
`define FPG_ODELAY_CALIB_BITSLIP_OFFSET 14
`define FPG_ODELAY_CALIB_BITSLIP 32'h0000c000
`define FPG_ODELAY_CALIB_EN_VTC_OFFSET 16
`define FPG_ODELAY_CALIB_EN_VTC 32'h00010000
`define FPG_ODELAY_CALIB_CAL_LATCH_OFFSET 17
`define FPG_ODELAY_CALIB_CAL_LATCH 32'h00020000
`define FPG_ODELAY_CALIB_TAPS_OFFSET 18
`define FPG_ODELAY_CALIB_TAPS 32'h07fc0000
