XlxV64EB    fa00    2470��}���Pw�(5ُ,V.�we�%K,�!=����3�o+�g�S���8�n!���A6o魂ǚ[$[�D!yY�Ω,�"7�f�t�{����b�|ouM4�@����ޯ��|^G{���U=��!"9̈���g?�X�2��bJә��*{R�!��"��*Y�|�0}O�5�lEz|?�h��N� #p�.:ʾ~0�8�������#F�0It���]�K��$�����
#�6ƦlJ� ycz�*��N��MS�j��|�S���=���:�)��^���N	^����z��MrZH�s����mI}��C�^�p�yL��h�0����8�h*��g^%�/���jc�JÛ�N�u��� 2������*�I�	#�Y	��w�>��<�D�}^\�O�Z���1I���ݶ4�#V��(=⛘H~�\ݬ���9s��?_�p�'�ّ#{i�=��R��k���v~��-���i�����J��]u�i%� ǟ�4�R�����e�(Vb����kT�P.E�3��� �O3�L�]�i��7���:��<��84_E_��]���3|�Ђ;��M;M�4�C��Fp&�E3��ȇV��x�$���m�C{ٳYˁ-a��4ܭ��)�V��z�(��U�%=��t���u~����Z�;��/,X/�8�%b�ȎO��� �@�&R <nM?l`G������`8�5��������X�=�$�GƢT���A�jʶ.��f��)Vt��Z�x=Did���Q�K��\E	)*��dœ5h���}������8%A�7��P�]�
m��ć��.wԁ����虛�`$�R g����F���ڬ�^���؇/bH�����Ο����aEg�*�(�,��V�ﵮ~౗��7���r?˽~�H��,��^��vo��M�G���}ku���F��쵹��Ym��L���i�����zky�'�)�/�nx� �G�n����tɂ��r0�;Eʈ���w�yaX�"3I��D����[��6�="Z�]~�&cA>��zY�����7#@�h�� ϥ��8)3\	���[w��L�P�;R}�>��
����U~//}��s�XmuB`0���0%Gf�=lr�ʈ݌�w����i*�����߰��ͪ}�5��׻G�>L���|&��3k�?}�/��Qs}�b�{�!i����T�����,.�u���np�p�B���@��ځZ3�r/�����~����b���T?����.���o2�sC��6K �9���Fm��q�/�� L+Ny�E�l�(��*A�i�f�p:?)-�9��(R���^�2� ���K�ZU�_����Mk9ך:��O�5,R�D�m���?CFme�$�U���D0��/]����s�j<-���4	5C���S)��u��.�,~�c#��.!���e7� l�PD<2X�<F`s��K��nq�Մa�HOO���gޔ�J���y�;/&�#��S��e��ջ۷v��u��k30A�Jf��!����`A������p�8��������;e��z:fi�\W��\�ĸ�:eV��ۻ�U$3�w��\��T�eGZ��EM��$eJm��(�9м�#<�$�Jn�A�BB����Ny��LQ�蜫Çw���{+��ύR͈�X�r�u(%�6D�2*�R�Gf'dz��q=��)�믤�X���r�/9PLQ���ߪ(K�B[�m�B�}�	�Ri2��@���{t�Ƌ=n��<�ֽ�z�F	��B]w�&����� mA�9R�e��'<�s96�Q�E]�ͬ������t9��2r��꼸��l��`�?瓥��g��j�T�Pۯ6�I�����j�ر��f����Y:�wg���1�����g�gX��4�n`��e=���HTY�L��F}?��^�H�&}>G�����j�y{�ts�F�g��~�]�_�u�WN�w\�RO74�Ֆf8�����mqPb�#5��MhZz�T�tZ4���D�0:F���>g@)�gr��e�*յ�c@���硎�1ֿ��3:�ZA��4wm(���|�m.r�a�O��%���5^h���\j����&�Ṱ�֍ɃEP����+���J�'
eL�NV>����o�̥��鬈���c(�7�9P˚&j�DqQ@����?OZ�\$�c�̮�<{5R\4��o��B�իS�O�P���H~�j�O�e�Z�������Cy��iwHÌ�|39�7��X8FA��C�������;e�J�?�ɷ�U0���s�S���,��jvm�r��~�TO�<�W#" *IS�����g���%R���mPQ��c�W,ܽ��ۗV���P{><�Zn���okF���'�h��x*^�y���Ub��t|���H��F\�8�����`��&���X�� '�̶yq	��V}i�+C y���7峽V�i�|o�Vϰ8�X1��]MP5z��VWS���2=���M��@K�I��꜓���>
XU�2���C�1���1�����{�o�C����������lx�vs��8Mn��@ni�Z�r��C[����`09K�d�]�*"Q&ĸ��"{.�5\jߘ��A���\�aǶ�y��_���O��}#t/�B� �y7��g�����U0Ў���yIow����r�����
���p�o�`w �5���=����Y�F7�B��s�Þ_�US�D���i��Vws��/����ឤ�Rs5{�jt��ѬG��1��Ul=k*ˆA�sEP�� �u}񓧽�-�
������$;Yh'.K)�p2_�5�H��v��,Tu�������{K�vo`�R�L����9F7���>(�ۉW�3��2hJh�3%!���w t�fl�u�=���EoD�f!��--	�����o7�����>�"b�s��f��3L޳�����%�߅y��'������b�{�	���"5��ɯ����nO�a0��2i庙��Q��HUU�	[���%f*�[/�c�-�������#�0�����W�U���o(�ʋm#T�+�d�<[�����5`ɮ%e�F����}{�S���^����[�;Y�Q �G�=5�#��[���8��`��f�q~RC�-W���w5�x硫��he��><�PM>z��J�üK'�"��c�bH�.N"F�8�H��sʹ<�L�͍B{	�"�b
1|Gs޾`HS#�&?�-��Ԓ�S�}O��:U
��y�B����Re����5m����qA�"m�~t%���7�'��`��uzY/|F�
4YϯP�7v�Qͺ+������K�+�����d�����*i*�_~X�8��swks5oeQ�d���y�$
�h�T�v�z9���.<����Lp0;�XL�3�$u�e�+a�?�Ft7�(����i`W�qt�VB$H�N81�tqe���=5����l(~<�+�pYeX�cIY�ܘ{
{�� �B%���'�k�J��XF��ش���Z�aLQ�8��Tn'`��͍��Z��pb��ǚ2�8��٢�Q$�_
�Ë®��)�%���.([~�ثo��\(���[9�(~X�38��ĜP�p��5�<�0�;>~����O��ń�cвqX;�/H�ٸ����ҽ8���}+���d��'X�w��G��,�w�.ċ@ŗ���dܳ��`�����r�wI���MՖ)��\fs�xr��É�����0�<�:cX�}9����*5����	(׾U�Xk�\%���t��mH�H��vL����~rU�2���w���A�WO�����9K��As	7]�j��W:��إ�4J�~�#���J:�Ue�<����?�8�vi|�0���4��*�c	_�0�pu�� I�-,1�o���އ�ϨR�r���v%&`�ݹ��6TF����y�(s3��;Ex[
Y�ˢǠ��w����т#=�
h�l��V�8�Qjd}�k�dㆠB��1��V`O�(�ێvPq�/�}\�TQ���@p"��n��,2<:6��O��/�K7�>��j�M�C�\����:��hq�'A���A��30!,�����-��-��@B��",��i;��&�:�:�����o�����oCȱ��$�1���XV��-��C���Y�!�"��2�&�>�o�P,��"Aei͑a�̵��o@�c��_9p�Hh����q�g0D ~6��+���@
vz.�Q�b�CW��	
��BM�<�R?�n
K9��V#�X@�	0�r�q!�aI2�9ϭ��߬+� �W!>j�T�ʸ]��r0��,�DŅX��`L��=%��z����Ķr"�uˠq�	�q*W49e{����&��Rs�B+��#I�' �1l�	��r��Z����*C����5=�*���z�V�ML%a-���c?6�\o�s�8�̈����PsH�W��O��舴b�^P���z=��e�k�z{���0�;����>�B����l���ܵ7�'�֞m�|�X�ؑ�\��޻��a�`$r���(�isj%�'����qty�i 1�l��t�\���#r��������yӢҖ`���\�R��د�$� &�����$��%�{�g�]��$�+����Rn	���A�s�j��az�O�����;V4fU��)���0�riuJ���T��r�D9JM��ZJL̂��,خ{f&x�<���#h�w	�qô�j¼SSLC>�s��<%�+P�7�=M����^���j/6G�g���1x��Hw��
Nbz7΋�d�x�$]Z����9�c2���X��9�&��;�=F-^�k=�`h��`"q�0Y�JF=�8�6�G��w�fȃ�QRo����
�v��!�d���ws�NV�#����j��桹-!4�^wq�c�t-�A����վ�y 5L�+K��RgiMv4��x�L-���g;6���w�sG�A� �A�l�Ep�O�)rk�N�J+ʅY�;7�� �Io6�� U���b�wN0-�D?�#u�D��E�ш�eV<�V���/Q>��}�,�k�˯�/���_8�5w�S���m�,�@�Q$`���i�/�5�갰<gå�~&��������٘��#q\�G�'�\�����I���Ch\�U���u@	��\��j�n��S
��i���غ�J9��L�C�gڙ�'c���G��p�f%�� ����.t��4#l�_��$�G�A�ב�C�Ę����#dn��i�tT>=h#��^#s�%��ÄTX4��]���27Ʀw��ͧ�=��']t�3A�i1z���G��,>ё�b0��f�'��`��I%�U:}�S�E���_
�_���s�v�C7�ȔuA��12T��RӘ�p�
0Ql&�����h�E���N�����(�:�;K�����S���
��E���;�e�����+�R�b��ȔT<�~����L3��cW�є�F���u�Uo�o7��lR7}�pdp��\M6��I\��<��|���#���:�۶��Y����:�������u�;��G�=b�,|�!{mg��&���E�z!S�D\ �]+/=cfs���e��D�t��/6Ef�b;�X�~�4`]M�eZ������͋%ۺ��?��BZ�:�I1���\�WbG��������Z���4�;T������OΒ_+�c1S�����F�>�=&O9�gW�W�G����OK���$[�K��sv��5�'`�vv�f�sS�خ~����t��K�
1������7Y�2����VYZaQ��=�L��Q"t����BV8�C`X�G�:�g_H��ī�(��~�1���p�y�j��j�W{�-In�ï�f�%D�|�Db�Y���ӥ%9yG�ݬ�׻[�	�R'�I���5u~����p����s��g�J�o5�go���-{a�i,��I؟�f�knݜ�I��s����<}�!�D&}�#���D�Քޠ�P�\����k��e��	5 �f�f���%Iޒ6{l���4-z��-$N�K���~ˑM���*��nk��Yu�ў��I�P��������-l�:�UpG�l����#����b���z��1hT�	���{w�~)&�O  41��h�x�H@Ǯa�r�����5�b��q0��9�8�yQ���#��1����ۢ�n<E�*�����"��1��%�ܗ#zX��^�gy���wMx8� ��R�TN����$D��1�M锼�(�j�ǫ���~-~���Q,W�Q��>K�9�:7F)Zm�ɝ�f�w�- ۄ���[��KB�a���P���|�ϪT��~Hk`�
5+�������/m*�ǘ�=���#���P�|Gة/�%��@�zJ�����H��nV����-vU���r�"Y�m(��s�i<���Mbg�:�!��cœc�7i�l�����V�'8o����q�z(T��'(<��@0�I���<c�P�Sf]��R	��`��W[��Y��o��EX����G�:��M�U�SӒ�;��d`�[�I��Щ�-`,]��<h��i��>2���������ahq�� �jyU~�p�T�v�W��V�bn=���
���Ģ]��
���!��� �]���Ƞf�_��)�RV
������#�y�W�e��ժ��uPt������+f@��,,� � Zyo�`���G�7�Q�Ǖ�wi�,m�٥b����;��!�x����(�v�"_�����^�-����4���^��fv%����i�4�����Nֿ�yۺ� ����ɸZ۲#`w�)Z�������ÁC�����@Æ����0�K�A3⵹�����c��o5�d��WF��bV�2̵�y�ߘ5���Y#�+�ٮ��.���a�~x��&O�������c밧#�{��Q����� mE; �D�̂?�����o�*��p�pɪ��L�J�9<|��ѧ_��`�I.�7�
2�f���7�#��e	S�u�((��bױ��ӹ�_ȧ�+�?�Va����o^@�(��<,`#�zN ����t�>Mm�X��ݦ��%EFt�4��)/4َR`,}�b׺*(��D>ӷRbLm���k445�Co`�dH"s��R,����@��L~�Z�r{�%h�}��@"Y{K�;�X$����㕜d���{�dB'��[�q6�O�^R�͖d4# ff&����G<L�Sdļ��P,"!@�����:��镸��oǊ����?�_h��ԧ�t� {`FBn�)��%�#�{��:8@!��rX@��FY���0�.��\�5�݊�m���<�OO�g�N�7\�{ �R�##��naw*��\�\0cQm8�BL�a4~v�\j�WS0���Ŝһê��[�6�rɫѢ�9���=�(�a�+��mjKŮ2<pﾃ`�7�	wA�xE$��=��{{�~!?B]�+S'��Ӓ�]�ҽ�^�����+7�Gb.|�CCwi��:տzk��bZS��h.L4X�$5R�$#wt:�pT�-��9׷�����ڪ��Eͪ���a��i`Uýx�0ӓ[�x!A\۰#�^�@��̵d��T���f��rq.݋V�D��dgҢ��ﮏB���V���:��#�ٍ�8�"n��aPE���A��g�,�	m�m�e /[����1)�(]�W#�Gk�(u\��A���V�'�6��b6���_�ٱ�l�r���^�;�2�K�e�=���wFϩV'��MWN�T/xV�Ք�s^b���  Uc�e���ϫ��\��aA���rw�AH�5 �}����#�i�a�}Yi1�g�]��@��-��5C-'vD�T��=*L�vh��J��-8���A��L���׶W*�#5������ޓ̍�HD&n���٪��k	Z�k�$���p�� ��Bo'��ѧ��v"��-���R����*��uMg�wNցZ�^��`����%��S��q��2ؽ�ξ��rۙ�q��.%����y��u�2g�}}��7��&i(��Ӗ�B�sꀎ忧�5��U
��"qy�u�w�g�lF
�<�Rh١���b���OC6� �ͯ� V9\v�����*%P�*1���P������R��N3=	?T�6��IIE49�8�GH��%�K����*�`�>�kfL�0L ��e�9,�����O(�	*�X���]� *�FL�.��j6(������WU�Z~�����Ӻ����r!4�ż> �u{	�.��4�k\gX��%�^��[2?��/���{G���������H5���kSa�L���-�mX���r�>J*����	V�˼|��B}�_�V5f���kgI>�`Ǟ��5�o+*j.L��]�]����(���b%���Z�=ۣRK�Y�K�%�=�m�a�!Oq���"{�K�a�u�g�j�6x��ד���[�E!9tvk�8�#�iH5?��}��~��Qh�q�l�4�2TQ�3ӡ��]_Z�-Q�د1���;j̩��q�/T7]l����n���{>�mt��!(^�p�nkx�mX50Q㳦gXM�i%���di�&p�=�Zi/�4,�2#<�]/8ʕ�߁Zjj���ιL'�F����}���C�
V���@��O7ύ�U��]��X����K��聟��I"K�u�A'�:�����nY^="Q��_'wu���G P�t��1Twl�qU2���/��q� ��o@A1+�N��m��P�)�
�)B����q��7��
�c�&C��L��-��@y�w7��Ҷru�]��^��/�	L'��{)��e0��S`S��J�١��T6>�p��z��_���Js�F�ut�	���zn��;rx5�n���"����0�aW��T���k��к��i72�Q[�Θ傁]^/�F�qb�4i?��Wu1~�?V,�{nW�3��{o�9"��\����r��B������5�B��ޡ��?��=���0��%>1�[l ���t��?$�t:�i(�R'���ma3�)]������}a%�����Tn�K��WS�Lԋ��\/��\�3.&yty��TԦ�_-و�;�����~�n���j͔!�XlxV64EB    fa00    1b30�G������o�'�?5R����`�g��t���Wַw�ɺ�p2��0�� \���)����_$�� ��G��BOe0�b5
���� K�	�i����_�څ�갶�\c<� w�?u�":����[�)?%�=W�V��Gb`)T�b`L�%O+�$�J+@o�|-��Q��<����sB[����5E�h��ãY��`&�~kW��Q�چj�AY�f��:125NJ��^.,�:��iA��~Y!b.LJQC��)?1H�	���/���&��Rm�Ь��O���dj~�?���ƭ�gX��c�(������;�������4��s��e��%��V'N2���GTŏzv�~Q�����ũ0Ĥ5�v�������� ��:��jh�+�X�����ty����nO�̽���E�AH�\� �{�Ǖ��J[�*����}�p���6+F�t4��|uo��쏑lѮމ��2hک�fU�%L���~E����r(<:�����'�������֌@~Z}�-�A��i~([s��(gTS��9�7v@���/*u3>~WW]�jQYK���23�
n�\ǶKo�$櫓�����[�?��Gv*ISD��'�o�>�2ZSw��6_�|����
�N���{I�#�ܶ���v���W����cv܃
a?�jn�⡝�?���`n1�i����	Ỵ�Q�E1-�p0�k�х1+o;a4Kd=�����f����嚢��.}�I�
D���͑$��N�نO�!���UT��=�����N�mh���wq��=�wZ��d!�=!�����.A�(Qx���ɚ�僩��xJ�����M�t������djC��˛��s���,�>�q�'�%��r�T$��������!��?ctk�� ��D�H_��/���y��f�J$����X�G����&�k%嵣�O��C�{��t�JY����gF�C�Ԑ��'B���ET����������yʄ�d����g�M��sH�q;��X�MZ&��7�2�'_��,�m4� ��>�(l-ݹ�y�>��ݵn�$�](����9�R��x�����&�9cEYibl"�6������?jp�Y56�V֪t��������� �m7wE?�bm$���N Iw�=8�6:�4���5-z�u����֯v	z��L�-�3�2
� F��v�`aͩM������У���)�e2��3�1z�7��+���zPD��dp^�rA�i`��:K\�k9�=����}҃�a,��XL<�JSH9���`菨�@�l���۱Ei��}���ozl��_�P_�-�?)ΈD��,4�]��"�7MTPn��N�j�������ԃQN�N�Fϛz{���G��')ؓ,�(�<I�ٙ΀��l}y��&ЍV�,���^j(�87���;�Q�+lB>��Q�����_u�3�>�b��hl��lP1R�_�c�'�I�8��B�!בVؐ5\��`C���׹,�[L�S������KC�#�1IC�n;�#��8+
u6O�{�g�zڂ	#ț8��+��0 ����_M���W�$���aH�9�+Aa�>��Q��'�_��2Qc�f���&��M[�P2��*�ݝ����XSUG�%�vM��B^���J�n��X���h�t�=\�=!�z�O_�{�f�@�>m���X�%�"�Rn��N���f5�fhk��gkk �rF�dmQԗ�e��5t�߀w�g�%V� Wɻ��P)z��գ}�:b|�ꛞ�k��}��]��wuS���Z� c����o��ݢ��'Ċ
��̽X��7P�#(�>�6Z��ڡ鎂GdY�f�a3����puW�N/�WF9YJ1ʦ�O�lc�W�:_�ݍ�}��&�x����=ч0�����%[B���"�LB�'ťsO�;�S�JeY �8�H2(��4������W<��FF�D��H�L8�neBE���H�=2T�D��"UEq��;fi�1��l��)�ә$GXg=��ݭA�ZZˉ��ؕ�_l;�`ס_�$Ē=���`E��+� ����G����I�ʓ�����F �w�&]��uh���T/���f�*N�;K��E���zN��;΅_��YX>�ҩ�3�~T�)�Ek�H� Cټ�yQ	<�w=?}�?�D���n�&8�]�0��E�������%Q���zA�ᗅ�]]=g����;d��'��j��LV.b1���.��DE�Q��k�칓��F�����> �����ItWnO�XH��?��V�I��C�L���2�Ⱦ���3�����T�-�A�F2��ZT&�&�jIk����N�E+O�ֱ.#)���&)0뼖7/g��\\��RlM�ZvJn@�"Yɔ�h?P�F۱P|ǃc~�.s>%8���� ���e�x����@c�ɝ	�2R;-,�f5���q��r��k���·s�&i��62�2x���>-X�����ؚ/f��@Y�c0�@����Z�Ui�7>U�����>s^Z����t����k�Ϳ���
i�P�ݜ߯� �k� 5�M�-�;|h�n@�!��^��t�)%~@=��X�mn���_]� ���'"�Z_�}= �(X�<m�6d�6)�ίn��H�^|1T7r�����,%~��獊�>��癋�| ��Ue�f���37.�=�� ���Ƈ��!�XI�ŧ!��$���h��5�1D����5	����=�Qn�2��3�2��G����k|ٞ]h���C�b��Sdmv�u#REH��A,�?RW�t/
����m6�+f޼ׅA�k��e~��08������R�+׼y�j�y/�1lLƵv�x�<DH�e�z"h��Ƥ���!�( M@����c� U�����F�R]	*��|ϹM��r��u���sVS�{\ ۘ��G�5Y�4sZ��%�)䤳�7*���x3��>�},��YWW���f�1����_<h�&S�؛Q[uWY����o�O�GE]D�-w�t�����e��w1��!(D��X�&SGI�����[+���8G�sez�Y����!��)�^8�ǋ�0�nl��[�ʶIʔz<�e��$��9�&-��-B^��Q�j'v\^�(5�TM�"+t���z�FF�)���p���frs�C}%r�FH��K�y	U��\��٨�4�ē�G�1�jSaD�J=�<ZU-��w�/��5�}���pD��35��s�������ՋZ�o�O	g�U�3���岟���E��΢�C@/߮2�����gQ���pڣ@�YYΐ������co(8�*HK�@
������H����F<�M�8�p��g�°/����^�4���쿎fZ��Ԃ��+g����]\6dhP3#6����O"f�7C7���WѠve��������(g���ݽ�%.M�������%�u���N*v��ɺ��9�*�L��aP��;{���{iĜb�,�m�2��\���$�u9�mk-3���Ej���P<c���˻这�M*Y�Z��3�� ���3��w�:����EU� 㔦�tK$8��v`̦�$�������VH��� ��[��3Y�
����	7@^�&���(�ߍ�.̊5�S�T�T3��5�EU���d|Lw �,�t��
����K�S�e (�(}�0�lTt{g��[��
:J@߯���+L9��޵匡<�گ�tx����F�Ep��Q��ɗF��s`�X���MI��7|[Y�.�筋�X�|Sv�o��������|ҵ�y��~�I ۝O.=���T�Wj�Ӂ4�m�;�b]��)[�f�\��'������ܦ^�,H\�G���t\�x{ۣ����_f;dt�����p�YID�* ����Ao6)8��hL&|��lp�[���
�>��;���5�6�@����h��d|t�+�_c?���R��%ꗷ-�f.��#���Ϩ�L ͷH�TƳv7��M�T*UuL���*;�K�w*��oƭ����m�Il�o����V�{�=8D��Ŕ�7�V�j~���wS�Ke�2��p�ڕ������\t�և����G"�06G��\��	�RN� �˙����I#�7��FB�ے�IuAj�c�h�c ��/��{�2�5	k���i����W��B�s�2�u��L�Y��i:�-�>	u�8����O���X3��5�#.`Nx[�V�@\]��������1�@��&Yn�i��=��VM�B�*��wL��ep�0��� T;(��IJ?$��C�E*�/.SR�����uGn�:~��w�D��)�'�,��іt�m"V��uQIݣHd������t��o�4��3L��gW�ԇ�Hj��uC��\!��^C�Ǚ�[�����P�
/%�6SY��-7g�X3d����^Q���xE;t�n�FX��܅2Mc��(9,H^=�b���E-H�pMǌR��B���"8ʣ_�H;�=�⚦u��9��s]U�S6��#Pv��h,<�qDR�����_!�:�?����=ċ��2Kt�`�.9�U���Ŗ�q3q[��C]@6 �Ssq0����s���F��+�+�+�!������\��I������ʚ}�^-���f�2UǤ�����pF�Kѽ�����iR�>**k]�h��F'�}}�SR������J�H^M823P�������X�:
�e��9��d�	���iO� �!�FGS�B�x0�73�iZNE;�,;� ��cI�CUq����1����q�!���/#U���Z�� =�k�Ƽ��0�A��3�[������b&�G6,S�v.���P��Q�E�dyZI����*��h����h��]2}6�ѽ�q�A��1�s�<S']�1�}�@v� {�,#>%��ɛ��+�����2e�toH�ʵ>�*�hI��j9fY�wziP�2Ѧ���J��{�x��S_���O[�@���\U<�j𖼻y��8/����ޅ�z����o%9�z��X}���E��DO��6d����a��\}#H�j�ac3�.9�Q7D�u�xp���Uj�o�J5 ڷ����8��@��h�k��;��/���^��-��K�b���i�j4Um��0%p^�����Cw$V����6�r�q��{����%]�����3UÕШ��JUl|�t�b!����bYVF,6-�R=�3u��ͱ��@���V�u�aXg%.p��h�xo�Ű����=����r��97XlZ\%�ɘ�O����!k�-����b��zJ� �p��t4�|م5�T w'���i���XEW$���\ ��]�Sb�n	�t��i�`2��w(������V���0�m�N!D��)�b.OF�H�^����ĿQ��z�j��,�5��ٵug����-o��~�g�7�F�8o�-?3��ys#�p�1=��E`{0)� ]�Wl�v6���*/��
,�?��jm;��(TF��;Ƀf�l���ʧޥD��u��j��4i0�Y6���45zioN�P�C\Sq�ò��]f���?�H(��%�����]\+-�ng���Կ���NX1*To ���A��:��0U�"�a��� ���x�خ��9}�~���HI�Ô�_a��F�WK1 BMO����L�lL8�VH�g�ri�0�g;��J�/���Lu�}]���xx�ig������v�����*I��� �T�o=Y�����eSԹ�6�E2�;���C���ԇ��ej�AYN��^�-�L?�L� X"��
I0�����a�N��5sj�P_Oe��j�˲�Pb�S�#L�w#�H���qҬr�����^N#Ju��QyKwt�+ً@H8��O��k���9��7Y2��F��O��v������u�,#/��� �$����[���u�����Ga1�sQ�_8k�*�u��}uGe�c���}���u�ii��f�P������E,W-q��jc�y�}�)�H����?��N�6�b
S�AlhY�[��w>+���qr�B#�-|��P�GK����֑���֪�%ǹ�[�:�W9�#�`�L3�N1%L�/�r��5��AX"�I)^y�\���C��������m���]��Q%�K>�x��&@R<Tx����N"�b�[YH%�����������ƶ��э�S��ރ���L�Ne�N�[�K���h�q�Q��kciqt�F���������-Y�c�����p�\$FU(�6����{�����9����waL��������tk��ϰ߆�ٷ������Cj�w�W�KA[��ܖc;s�O���9�-w��R,�.�t�@���JF`jg81��1�ų�2���.ك6�1@�4͗-���T":dj����C����h�U:��2�e�3�J�X�FC������3b��x���Bn����6%wUu/��!`<'�o	R�.���2��*���Y!dK�"�����h�4&���>����z iz�?Q| �`�@3�+ '훟y�[_9q����x��̅oK{>��^e���O��Q�H�C`��ے��ЫuZx�3���J�ˌ�}�zl�W_�͉܃�ҋ���>����"��_�_��=���C.jGs��0�n]��0�0��>K��E/	��h���OWy���U��q�Lإ13f��Џe�,�R} e[ǯ���v��vVD����_�ixi[�Y"��!P�y�R�vxĴ@�[Y��󙒠�Ϸ�3��(�[��������׮=%θOmɚ��. n,��_s��r�K��T9�fDdIې�]��톤�B�~�Y�<�)QG��1T�XlxV64EB    fa00    1950G�H�w��zG�&ë���\� ,�(aea��!jy�"��K<��JC�u���ZE���,=\�Y}�pv1�t��b,�� ��|b_�6�5!�C����!8�AQk ��3+KR�[;��KQr�Q�l#:&��m�sG���O<��������G}�k��L��@�o-�˵׾'k�S˼#���3\��%Z�-� ���$�a{�%ZB�� {�O`>ⵧ�b4�a}/yـ���r�������)X���co3���i���Iow%U�9R��ϭDMW�ӽ>�g��zq��N�Q:+:���)���W�����;�x���-yh<��R��s%v�'\3����,R�s|�5���'F)��R�wM0�.���o���OhA��c=�#o7����O��R}���
���քh/�>��&��ͺ�3�I6^Ջi�J��Ւ���U�_Cj���m�=�p��������p���("O� �HW�k�иu
�O�[�w�;�γ�<���mpL�Z}v��1��J�����^�yS�bn��7~�d"���W�M�Q@�0����ða9u<ħ9��7��b�50$�fI�3h쟯�ޤ����-�ɍ�i�<�L 2NZ�#�n�Z�"Y��z�Ȕ���+����f߄�+7��x,�H�	eY�"����'��תA�à`; ��2�����}���R�T�)��v��x1�+T`��pj��D�>�6bc��&]7��rL��{a������P,L�K����@0���|���>c>����H��?�H[|���Du'�Z�l�쵴�4M�7g�Fn��w^D�Ef�ʘ��P�LR����t���R0����g����_+P��2ӕm�<b�』�`'�ɍ٬~T�O�x���tk��ɚY�>��J%�˿?����_4vO�u�K�D(=����`j��1���]h�����$X0W�I\T*�S��g�Cb���[�Z��0ӈy�����P�H��	�ߜi����4���l��� �(���~��֚w�.`� ��BQ������AC �	1�"l)2sJ�֠Q��d�^*�=BK��$�~'����P4�8x��ȭsĈ���/\����1�v8"�¼.+l d���W�e����)U,�Ձc_G���)�[�?��<���Q��[_T)}t���e�A� �)�o����y�j-��q�UL"��qat&B�כ�{jB���~x�^<9P�%�ڢK�p�I��(xM_�T6���a�brP/	�8����75a�w2����	H?�q��\Aʪ)[�e����߭��*R0x\�"���T��)��Ȟ`HtؚEm��~�f�Д.Ik�q#Y�p�8y��L�s7��9��H,�ͭDvwCɵ)(�-��!�m?W�K�%^z2�y��ו�2(�q��Ԝ�a,��B�ƴ�oҶ�`g�;8e���1�eЙk�e�D"�o�'��3������#z��W���:+����b���?��Q�^Q�#g�D�!z��2j�R~��*�>!��1�4��Z�D�ü��)��B�aE+~3�X�-��Q ���_�g�Z,yh�(��=�p(wad��͋�q3���b��
��T�2h`;Y����|����NkD�Α�������T�ͳ)�]�;�����8 hԧ�A��8�6�,l��e��}ӷ��69`"T��׆;˃�登�H�u_���|C�-)����]ehpX�o����¸'�K�l�J�E�ۋ���'|�/�+ե�x���]�`]���ŌY���A��@oT*� ���;[^�5�JA���p����f������:���	@�99K*Qx�� 9
Sk���"������>��f�R���%��!�!T�84]�uw:��D>�m��))/�~���Xʲ�y�bw�[�U���o[ѿ��ڱ������S�� Q���VA�Ue��W�`��&�7G�� ��mtEu>5]Kd� CZ�L��0�}΍|ɲ��'������9ج�![z�+�S��1paU�Q�S�Fl7 �,w j�7�g�΁��*���5�pK�f�C33niU+���O��+�ʪ-�lhp�׃0�$IJa�F�?"
��ޢ���zK�e��d���53Z�\w��w�T_Qa�ֳ�[:��a'���eM�O��aI�R��FQ�C%�|0:�Id���P@�7� 7A��z������.	0=j�m~n�N��h���-��\��,Ɠ!� ũ���M���Cؽ@��?}c�в��0Ag���=Lߕ�c1iy�O��]w��}a���.���1R��C^s|=�>�|$޽S'Z�2��Pu��<o�϶Q�q���v��ƾ�5p�+p_�QM�|�C��u:�5�*2�M���[6#���ףN����z��J~ ������v"6)$jޭ������ DU=J�̥���rɸz]���_� DA2
/K"��a�����?��x�1�A̅�ؗ��o�b�/�Nr�wI�\\)���:H���7�\gJ�W���,}�(��JNQ����Ɲ])���?D��&׎D(�9?-rV�:W+ҙg�=$���|�Ĳ7���8Жw�����燐O~7��R�Z��񁸘0ꀰ(s� lӠr٣`�n*��a�:����A��I7 x���$������m�o	ٶ�,�m��R�kLd9�H����mc;�,�.,3K��`(#���e�u�q��W�*�1�m+��*ܨ��x|ނ�a]����y�|?x%3n�D�D��·:������)�[�(��)�ч��3j�r�@��ִ�����9��ܧ�8�K:v�-L�}P��Ï,}�fJ9���:f�ȧ�f[��M��kpc�`�/bb��D̏��P���}62��� 0��%��&��W��Ֆa��&�{��}��>)r��ߠ9z��Z�0�U��#P/D�D��2	QZ�N�Ba�A^�h_��3���r���I�:FAu��x��p]���M�❜O��N��YZ�AW�=�H�8~��8�2[ѝS`�����-\T�b	�����׾X��R Vw�|��-ř�1��bWƶ�}��5i�.�ւ�F{
l��֡�$��9�\����
6��J���B�h���r�8׏�-�-��Ř��ݭ}���:3L�S���j�LZ���%-@��b0�h6�����_�H�e���9�@|΢h�Q�8˼�"-������%���ji/A��6�ojdZ�������$&�|�A�+?Q����R_s�[*k����ꊃɫ�-ʝF�CaH���?���!��:t~��罡�jU�e{V�Y���w3c^o�N�Zf)��&�l�3ۈ/�# 7����8����Aԕ��e�_D��=p�m�hGx��T���~۸����4��� ��y����
õK-[��c�ƙn\b%�!��2\�7�|k����G���<�S�\G���.CҪ��� �&�ԉ!����n��Y���a�`�\�b#F�By�X�:�P 2�U'�Y�Zz�iY��R��a�P�*0�9z��$��Z�E3xP�B.>O���c���Zb��_�����-��r;*��Gq����]��"H��Q���Б�c�mP�2�N5��E��I�~��\�IE�8.�p�=}h��?���+E1L�� ��b�̎[>i����k��v]E��P׶��B���-��"V	����?
�r�d�.c)����Y��$(����^<�A� Xf��DEEfca���o��)����������0m�͆l(���H����N�)|BW��z���`�E���u����ݔ�[Kk}I���>-�����"u؂ez�M���9�������e$x��U��5��BŇnD}T�i�IK���G���O�߈H���r��c,��e	��%��mE�A�K�vY�NO��aB���̰b�����E M_t�g�'z�X���P��D�Og�[c�SǏW>��<��6Q�5ǦN��ؒm�sl�08�K���Z�NI���`j��YzM�[�����1��N���O�e��N@�ب x��Nd�Z�����7／1	_m�W�u���;-	��<#�b��u��dd%F0&<EJ(��Z����p����]5��HK�L����Ki���U�N��G�<�>֙b�UB��
7_W�����6�FŖc$�������X�С���K��7��[fAЙX�}�phLC
�7��@�B�#w���"�L�'�(�'ֶk=�<<�5�^�=��=k��-�w[(� U�����V��Ǖ����i�?�Ʋ���g��nm���sg�P(���2�*�k8���o�d�d�4Ql��W��A "�l"%u��n��'SPYwU6�$\�p�$���O���v�Xp��yJ�[�Bkv�w���?���*�oP�LN
'��ȯN���_�[�P�Cy�ye��p�۝?����K����a��j/�����	-�c�-�����;�E�v�-��1�xt6�P؝89��0�@R��1CK�ů�Oa�5	,�%�K�PrhJ3�&b�y�8��|�Yy�O��S���''�Z�Ğ�s��w��J�0d�y
�����h����?X`{�W���è�d$��$�(	Ԃe�8���ɊmK{D����}�|v�xG���n�pt�����r���E����X�*m��}�5�1��t�
��j�Wa�꣗4��}kRy�N����A: I�N�n|?ht�A��mߢ�֒y�⅕s�T+""E%�̍Tp6����e`��Ǝش�X�ί(�R�r���Ǭ�9~j/����0�/��U���x�*��=��K�_Z�����u'AlhLf�I83�����`a�D7k
�J������pZ���H�8(�����'r J4c����k��`�nL�݅`�6�O��/]]��J_��<�9���f�d�3�9��
�j<�o�@�o�T�T��63�4ǌ!�꣡�$<clܢ����1iu�z� �ZG��IY7�6b� I��B||Qq��>��ΰl�pWDؐ���_��,
#�C���<�hBw��ű (�K�?�`��,�ý�E��!��9??6%�qR����
��z�r�;�[7���m���ԋ�Yd�Q���r0�=�o�&�	�T�/�8�(6e$νK�ň
5���?<56Gx<�S�֡Z�{dؙ}�"�+��>�����{|��у�ۄ.1B���~X�a �ЂN�>�U.s��B�*���e�/o��_�
yQ�?:��
\=+����0r�Q��,�񍺼��E���[NZ�>R��	�~`R��e�9P��3�2O#���d��9}9�i���:���~܅e�m@? Koe�YN��C�ހ��=��%�g�z�G�)��z�!An��u0-�<������gy1�.b��3�L���L�(q��Zs(���wV��ɞ��؍kCS�c�z�0��/=����e�Q�G��;ˀr���V�{s���R��	��rȊ|E�^`e�;��Q��R�m�h�G� ��ry��m����Cc.;�K������zm5C����?��J�ԩ���%c����*�e��҆���t��@R���IkN}���bLGXt�a�^It"��x(�IةBR��jX��-|&'�Tm^Ľ�c	��*�O����l���n�@�ʒi�-���qV�"=�&ҡ�%�q����I��T ����~��U �<⶞�b,mq�"V�ǐ�s����Lc��t	w}Оf�
s%�3�A�π��=@�!��[�'(���:��X$�=r$4N���3n�i���y��y�$��:H���f_J6�*�)E3�y"׮
����j<�`��"`���w�F]� &�	G�
�|8b���8Q�9}�O��Q[��i�ٰ=���8���g�^v_���E��_ü�nS�ff~���:szivcLC�~��˳�'��8�;qM���;ҭ)ص^$b><�����c���4;�,�,qD�
��N���=c�	F´Γ�s��kB�W��3� ���i��<Oj������nM-_}ۣ���h,�]g����,)6L׺�j{���� � ����b��~��EmRpe�2��������RQ��B����Mu��v�����_���hz���ȷ_O|8�i�7�rW��{����W}ҏ�܇�Rb0�k��Ǉf��1���]$�V;=��y��}B�s䦹�]��\�L9��R\iH���Y¿A�B�:F0ǁO]jN�"��&��_D���"�z$C�bR���vҷ��$�A|Rd�֧�w�֚�
l�)�ƌ����k�` �O$�O#���Q�KB�'�U;�%�)��XlxV64EB    544e     ea0�lg�e:ࠒd:�(%=�0�M��]����ya�[&]�fzR�T�( ��f�f�q����Cʺ�-Q6��f�CŠz1O$��W{vf�N�-�N����%)���
�izR�!��3Nݩ���b��[e
:�w96�y���0׼iݹv�:Y$�bf���@X���p�>����8�6W���~H+��#�����DY�K{
�;��m��Z����1~h�U��cX���įŁ��`�No����k���A����"�����qy��&���|5�� =ѿ�
����ߪ������1;�/�{��v64�@{9����ӹY�f4�}��v��:�9�M����;z�����NU���w��TQ�*_�0[,_p,�x�	6T���d����x	Q�?�����zp>r�3w��JK�"u���A%L����	˩(>ڢ[�2"�X�����c6GUX)?Z,�[�w��z:�f����}�L�(L����v�Q:��w<�Y��rI �)^旺z��[O�3���9 �e��GwZ?|{�� ��߇  ����lO��+wf7c��y>A�\� �k��C~� �K��9S��8�;��|hG���u	~�s�������%îbA�vL/��.\���|C�]���x��BW�F�[G����0����ڜc�ll6�F���Վ����FqO����SO���<\����:o��4��~�|���ԯ��qhNv�{�j��ؿ֠���Kѳi�G��?��5��?q�Vc���I�x���i�H�Q�uB�}ާ����^��ZY�Yv�-�' ��/�!�1T	 �~ܠKa�}�B}��ɹ��x�*���L���ۮG8c3��Yn��?�
��E	N����V�����D�N$k����B��Il[�k��b�ap����R��=�dJ��G���1Dm������W�w2�$�_�t����l#�|��=O$�*wB�2����h�L��y���QهE��O�D���Х��FdW�S��Ö���Cy����6U�9Y!Q �l!�Q4n��eF�~�(��.�JE��@W:���'�ؼ�&��m��*:��e��	[h���YFs��	�"&�bv���Qm�f�ܕ l�)�U�R�#�ڞ.?��,�i���S�/6���K��|D��0�xQ�<��+o�_"x��,o�TEG��6o)�a���&����#!]���~}F:�N��C�V����a+崝1��Ԡ��:r`J��P���Vb�{��_x:~�[YisZ��F!'7���QҊ�4��a�\��m�-��֗�ڑR�y;�.ֺ��Z�~TS�D~��.�Q��5 ���%���E��*�
fk�_f9I������-I]��<�^��d�o��ϡ��)���غ���/��9�E�8d��k}m4_��.��n������m?�_e��ͺQ��M��p{��������b5� 1����L��=pF�NVWđ=6�b�����K�_7�㼩���ԅ��a<��s}�7�D��<&�`?O�]z6�+Kh�B���!�2�M���>������]��ɾ\p��e3˧�q}.�M�j���X��q`���Ft�KՙD:Q��6_V�Ov�Q'35l�|g�Q�F���A]���m��6������z܇��$�Cܛ��^������톦�{q8k_eY�*5���n츑gxu4��}f�A�W	K5Y
�#�a2�O��#�?_p?}+�@&}��C����-f�؜^a!�/�����Lqn�-q}58x �E�D�j�Rw'|5S���0	�0�_�R`&��^c��8� 3��ӫ��(������WRG����>,A�hW��7>6BR(ڒ"8 ����|��B�K!���֞������q|݇)��/�aSsz��7�O�� -�4:TlE�5�w�	�[Rb!Uo�KU)���N�KJ���hGb�gX�Z�Y V=��B�mN$C�{�����c]=c�����C		Z��?�o�'`M��⻜���&(h�)�{^� �S�:����3l�F�E�>�2CX�-{�~��+] |�3���>��6>rG��n�� r��"�Q�y�S����H��7����Ֆ��*z�'��p��B)r'ET��`�	�����)�/9�����5��5��
{.���#t�B��}e�Uĝ%m�VEhQ�תQ*J8!�J3�CP�CūͿ34@��N�e�(#ُ\��O���9F]��O%�)	��/o�΢!Fº�f�gEeC�䑙qzkw��}�ǎu�oi���nsq�=�Sϝ���wX���Soqu�cX�7����tI�5�SG3� �5<���ݦ���������'�������W�<��].3�&ߵjI��؉7e�w�R)�;Y�t���7q��P����n.	e��岻�Y\�ב>m�K��l���%S��:�/��")��b?>i#�$�~+�.���}�s4�_��+�=�Pu��rgw)OrM�3�~ҡ5	�Y�����M9��N�Qk�D�Ce�}��&=�-��?fiD��d��t�u{�����X��)B_�q���ײ�]a�Ĳ�^���AY�3C`�Px�� :���l�����#?��c<�f�B:_ik|��Su�s���|N�CY�h�������R���0*�0���(��xn���+a5â�O�"�����vtπ�Ӂ��?��^��0���1���96��q�B�u�<�{��@��=yx'�o�;��*>Hƺ�C��^^��i9�������M{F�S&<��ƎD-�}�� �kz!�!��tq@4�s/�&+(�hU��� �aڒ�A�*r�H�
&;!tSIPqV�mm�(���j��;�A��Q�q�ǁ˔�8bEr�$LH�ݞmt,T�d�׼~}�L�tx������R/�<(�FF`�������!^��쓒�b�Q�l�c�`n���0�U���J�TN����`���9����@����pi�%����y�ӛs��������6���A��=�M��T"��!���e�-#�Ȃ��r9��[Vꄡ�i:"�n@�,Y�f������?j_z�1=4�v��s�v�{�[+`Dp&���u~Y8�<ق�/;E�z��K��v���sJ���A�`{a�#R���u�ǎwW�b�]�]�sB��(�y�����*0^I�Ϗfub C��4�5��<�G�T�ZZ����i]���e�Z$����z�tm証�z���CkE�^���"
�-u�#(~=��uJ�<vxd �񽺕(Fϵ��c���١��m��R6A�`ե���]k�X��x(22wD?gB�IK�C'd=������e�h��{~�,��ѭ� ��`��B'�e��й"#���W���w�ױX�
�gtR9��Zk�7�	q/���t���Ƥ�9�˃Hb���@�����^�e�q��*����������%�;F�W*Ҏ�mg����z� u;�OR��e7Ej�ƌ�>�����bάP��u�gA��n��O(W���%ZT��!��~�q��wP�vNG��2�b�F�薵8!�I��ӎk[ �84��a���_�y;Ә��~��LYx��b�xS��7�%���0F�i�q4�Hnd��ze]�?�