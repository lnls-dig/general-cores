XlxV64EB    fa00    1790���^]M�>:w�tO��6fWN�
G�nh�d
�����ċ��y���)�1���li�7�MH�9o����F?Ϫ[^���^/Y:�檓�o�8̭ݙ%tڻ-,9�0j��~� �f4�cV���� �h!�u��V��NLG��^C�Դ�N}�����0B�@|�F,����Z&v�ŁB��Q�Z�Q/��v���� w���2eo͘��	���.�m���p����y��Q�Q�|t��R/��[�h���m�y���"r��|�}?
b����]㝝5箂�#ܩZ�/�jz&B!�����}g�I\s[Q��^�.ɟ��ء�mC�T�P�ʣOb6"���k�yy��^��Г
7��^,����59,�*m��
,���Z-�YnT�;?�v�H�fDp�x��LW+�-�r�f��vhB�����R]�z���w2�Pu8s�S|�4��@��+!;���z���ܚnu��:2�}��ؗ�Cn�I�K���M 6Q_$��JR:v���>tN��K��|�-����N}��1�$��*yۂ�3���ץ�'r��Z��и�o��J0N�e����_g�h��y1�z� 5�%�p&��6�L��6@�]�y5�a��A��)LAb8� mtIM��!r-�sM�K�y�l� ���~�+w|�](� l������0O,}�4�E{v��D���¸KS����I�ED3��#���#O���"G^
%���T5���$U�e1����T�Se��ua���
��T)��n]��iS��G�y�Qv&ɕb�k��d:O4L,�q�$ɑ$���!���J&��@�#I�纮ϴa�(����.� �w��r�QCg�� Lz�'��[�S���STu2�;<�zR=(}�:�g��<��R!�"����9��F�)�+M�e�DP�rN���g~���ϋ�&%����cF�TDA�%)�?cv�au�<[�}�F.#����o���A��[=}�FѴ1�!z���-4�O?���͏�f�@JJ����2�Wk�t�q��O�u�����{�����e`��=���X<w��u�]�+vh�χ��
�Y>u��z/���Uwʴd��]*���G�[<G�[y�B�����1��@ߥT���a'���)P�}Ik��}<����bv�-��#��&KU�se�3(4\��.���b7���P�
#��ٸ�i�\ODf�k j'��a=*�[b$���v�-9�@�/v�dA��Oo�3Sjwa
�٦�=J��4]U����Wؑ�>�1T��� �ޯVW^g����Y]�c$i	ݯ`���U�{����V���ׄ+��ꨌ"�*�Ur���ch[Ƭ��Q[M@�n��x'��=+�Syq̍��m��V�k2ݭC"�2���"�;o����`�#��~1�z���^��966���u����x�b
�n��d�)]F�q�-�	Bovi�����P�`$��]0��k�T��ZlAߜJÜ�St�;R�i$�$)����:.5x�q+W����S2h*�w)~���ũ�����:�lW�sK�c
!�؂�s��S�H��yp��W�#�6�]�G�jNy%�"��K&��' `ĠP>��3��q��RC1锸I~eg?���R��x�����Ͳ����+h�eV|&��d�?�L7�ַ���ȾAAT+ 4H�2�TH3��q�����p|�,�:�%Q��U����`�]x�G�;*��!x���XL�i�= �4���0�,������D�$%.�+&���U����C�G�"�}]n��4��/����0��˯�#�?�۵VE���9�,���]nd�7Đ�>f@	h�7	|c*�Vàc���+�!F�3��$ߔ��A�1��A픗�)!�Ls`_��Zq�|)�:`���|������H_(���^B���9s��7���n��KU��KaU�NK��ȿ��#3���G�{o[Hu�hN|�i��׸%?'P[cH~�8�3�W_���b�?�X Q���}�d�?A��a{HHM���}.Ȑ<��4���f�ܹ����a^8����Z����, 3_4���4�Jq{O-��5Ñ�	�M��w���K(F�o{.E�[����4�׀��>/VN4����sђԭ�VO�*r*�C������s��A�Xk���:��LvN	q�@�4[5��Y aYll,b5���C[���� �='���a��=;��-��ş�s�ޱ9��?�2�B��$��;�:�+�eF^�盟�(�	b'ń˖;�'[�b����e��G��tG��s��>B�b����Y��"����B�t�H�9y��$h|i�"E���}�f�i��K���I��<!�|��SqC�?�ӿa)}ъ��)\�(�C}_�gJ�hX$�%�q�zsR�(Q�֎gu` ���Ě`Ջ�"0YCzg�,��[�خ<�G�w2�۔l���u K5���%�28���t| P.|�G8s-��c��oS�l�Qf18��4�5�C�(7�^��Z�bl�g�}o�O$\��oIpI�r3�B?>���g�W�c���y�"�V]
������ER�O���O��'@�@=�A�V�,�-E�&������:0ҡI��[h1j�P�ٺ}����]����]���l�X�w����q��DxR���\���Zu9���ҁ\��2�������~�I��{�z����2��S�>�kYy��^r�Kp�uE��z��L(6�� ��D7�(v1+��5/���tr�N�r��w�[�������^�a��\/#O3ͷ��S%��q�"��{�h��Ʂ�9\ip�[6�9-�Ҭ��k�'��vP4-�mVoNtJ6'"g劰:��ԭX����%�uR�ޱ�d��l��	X�x隄<w��I�l9l�M_�(�D�e�ש=���~Y�s&[dMŐ)1_PI
�3C��5�b2}�ƅ�U1d�:*n�(Hj��b���c�ѷL��[�o�6��3;Y�LN�Umf�q�kHɎ������B7�f�^�.ov`�b��q#��}n<�kYH����PZ�|���Z��.��:G��2䟱Ur��gD]6��	�H�'_�����n����Rr����ޣ���\���,(�*8��_A��F ����,��"<�~h8� ��ͅ�2R�S�U��. �
k��W���1{�TEב����\ O��zPȴF�����
���@�[;X������[}����Z4��h�����C����0r�F�`�1�H2I�*�U��_���0`B�>�Af�&���
QB�.���A91n==���lt�0���X!6IN ��A2{�s�6�e�>K����*-vz�i�rδ,�3c˺�������������.��i�4�����_*K�]@c޶�¸z�n��7oL�-ȱa����&���H�&i�B!�t����q�1!���``:���]R����=A�!������f/Q�f��)e$*<vB��_!ȿNy-v�����m�$�<��\�P�5��� #�\qP��y6�Ö~��
���3c�`D )oFS�P'|2åN�2:Mh/���:���+]	�����l��^�������� ����#P��v_\"\��q�}����St0��HJ�ת�hw���'a�_�^�	����Ya �d���g=d��J��,j�M�	O{ߞ�Ī��,Kۓ��>cNh"��<�S���G#�6E�.��ꬽehVT5���R�Ѯ2%����շ��{���fG=��I��=S�(�����µ�As��,�:��񡞦�lo�T ��il�%�̲�"mQ��y�ph	-Pb^@��MS��{r��,5����(^��=R)ڏ�Ŝ1�'|��)`�R��h�G��a��v�)U���
)�i��Wa/�����}_ܵ����������7
�a7y��{n�:�W�rS��I9u�N��� ʼ8�p�Ң}�m�r�O�L|aV���`�+P�zȆ����1�C���M�	�5Ð���H��r7�r�NU�	��T��|�gtB�Ɏ�6�PJ�L���=ɠ���J)���Q���2�G�r�4?s�9�ua/��}+��E�!��BC>�a3�� ˮ �7i�RB��%�Si(��Azm�h�?����|���A������r�Y�]���N���j�	���0T�1��l6�$f��r-.��+	�e����Wl�H���B���p��G��ekP
��g.�o ��εb{jGh@��"�����/W�~?}��X���h#~f�/~f����hr|��/i�Z�=�$��.��6&8!�%b#�)�g�@!T.u���=�뫥0Ǉrb����V���T���jMP��in2�Yt�����Ѩ�;n��[hE�C����H�J��F3J\s�R�o)K���5Կ�R�	�r��跀��Ăn$h3�:}�j�����*������A�T�!S�m��G;���NM�\7 Y��L���9� c�
)�=�֯�X�H���0{��
�[7щ�@�(�C�����V⦶�א�t��D��/߽�q��&x��=���u^}|����B������l�á�Rd�$ ����xx_��N��yF�@5/���˰&�.�ыj����{"v
`�A�Q5�A��;���,��A֣�%l7Y��\=��7G�RWm	���4���V�I.�� �������OݚB?\�~��u��~2� �]�b^S>z	3k�S��Zn^��KƦvc0gU��k�4��`�u��)0���gA>#�s�14�:$ʃ����b!謺���r�����0mڂŐf T����RᏀ�x�kJ����}�D��Ў��4��I>\=��W�Yv�OZ"6$�(�o���d���������;�Lz� !Q���Awr,��n�KH�2 �,S�1>�x�-�I�.~����$���`��G�t��"�gk?NV�e��P5/g�J@��nR�}�R�`]'�V������+�iU�-q�_�U���H�� �qw,�z��ԓ��`�ե����#�(�	"��N@�ޕ!���L���5�l��mo��\c\8��H���n1�C��6�fK@(Wd5��B>6!7�y{��9�A~o;�����ę���+qp�H��	_�����XS}ZJD{�Z�_1X%@u#c��YB�.�dM�.�o����ZW�H����j�2�X�����މ�")@��ңLr��j�'�iu爭���Wh��\���L{���vY-��"�m�E,�k%�H� �/H�r��5��1��I����i���@��H���D��AM.��%�'*������OV<5���@�/���d|"?M[�₅�r�l<�/���2�����&����~��^$���_���ypU��g��q�X�O�o3�e"�ÆRU�G�������.������cǮ]�v���8��B��`�]7ŀi{y}�B8����Yc�#8+!�����`���Uȷ�C������<�A5���a]�t�}��z��j��ƃ
�*q��3��d�aV�k�"�D� ܥr T�i���쉳/��� ��*�!C�+���by"���C	WuX𚝞ݖ�ѵ���7��Y��?Q$�LS���Log!;ȏ���b�6O��DՉ�]!�p��IT0�%��P<=���ַ��M�����������=�;�1������
2�D6��E� N�����D]��Q̀�1
�j��y��7�Ϡ�C�K�_#��h�-2�`q{B�}�N��6܃a�n%0�G}����;�JX������챂2`7�s�/�~�᳌1j~����kG���^��t���om�8�2&���ن���^S^8��򩁝�Yk������y�x�y! �y1?`~ܘØ�z�&6XlxV64EB    fa00     5d0AE~�5?��E�jFL�8\���UO�C��zʋC�ˏaH	Z{m�̪s�{�A�:�U�:u���91އP��df����i�s��\��ا�4^S��ʜO����������������jg���I�QV�RGN�l�	���a��±]�I����6��2I��;�@}?LF�I���
q��9f���;�1b�>:��5��_dT�Ӄ���v%��+��1��t��3B�a�,�[���9���r��(�2��I���/'H�Q��mq�!�1��J��,���y�5g������Y��u�j�ݠ�1NW���`W*�ٮy�����6��L�6���`��!�}�S���%.$��l�'Q;�`�n�z4BQ�u.🛰Lj5��|�j��&�bA�.��g
�߀�����⨚����dj�)�fj�z���uR4�3���=�e	W-/"8������y����`��rA��b���H�+��U7� M}T�'5��|GD�������"\ɯE��I�Hy�IF�1�5s�0���o���%���>����W*��t�䌥�t�;�*x��q j�Q��ƭ���zd�:[�͸��oJK v4)�Qd�$.��!6��=�\�L���ӌae�	0%��mbLM���`TD3k!T��·�YB޾�z��rݗĳ�Ky>�{i�3�;Jz�2�n/�*�ӳ���B'��b� �v�ez�<A�a�V�$ȉ����Uۉ1ʃCS:@(�B�(�J��0�r߽T"���g�w���6_����B�)G����6�"k��:(�k8pE"���7389g����@�`�+�������į5:
�X��,��	Щb�j�Ǫ6���`%�qsӣ�]h����������>�/�(��@r5�b�� �+6.��yc���8�k����'���&]�����V>}Ac]��|�a=�I��]��!8+\+�o�(u�0�V�0�#g'���ؚJ!�ZKE�,�%��rA�s���~jy��H�è�p�{��u����y�ˮv�;^��TBp�6�����U�!�tP{[/R���T�I�1��p��z��UMP$�0���Y����ʆ��+����{C*�{~��b�en��ӯ�j�2Y�;�xva�l�\���=t��@mZP�]
��۽n��n��]VKG�n�(u����;b��Z��;v��Wg<�o%znq��6R�4�H~�����P_IހU8N|�c��PF6�G�uOOǘi:�*_C��p;�&�زy��h_����p����	qxx5��^)�>
�r��Y�?;7-R�����z���z��g�){���߫�0;(��i�
a�ڐ�KEF�&�t/!��Kh�9/D�u�e��l�pL��Y߲�)�e�Z_�^�D�yA4��R�mj7�#��5c��:�`��0JtH�f(.Q�.Y{���wc������̉DAaXlxV64EB    fa00     640I*5���P�������d��%JO�ǺrBSP�eᗠ��,�6B�b�n\�0?��[)/�~r��a���	��<�ԬxMO�Ժ@�R��	��m)4��P.�Q�.�L��^~�;�ŨNhNV#]�/Bb6�����c��Em�`HT-j�G �D����ҫ�L��z�)t�����a��a;���/���c�S���b\��\~����״s����bX����9��mg%�PQ�2����)t�}�hSF��.����,����=�	%'�K�%��IݪP�H�1[����;킌��#�J%LΆ��tz�1؍b\�+id����X���Le̘��1�` p��^|ȗ����%�	Y�m�͠������<p.����T{�#��w	f�D� "���f��@Ð�@L̛�$]����;��5?ǵ��u]R�
a�;^e=�şQbӲ-��A^���W_i�lI��GTCail@�nT����a���ԦPY���X�#J��S�	���H��Z3��/t�땃��{��>�t����A#j进�5P"��ӻ�:ʉf>4Qd[�����I�` ��m����z��k.�����m}4�~�	�ĩd��\�2T�8+3���"��Ե�u̴o��wڷ�[wL-����F�(o�H��{_F��*�^2���>>s�f�f�v�lkC��0�G�!8����_�hf&�C��0�u�e�|���p��M�|^����T�(�4����`3ek�H�#=����ލ`��厦+'�NT|���~��J^�냵�p������r��Rh����^�%XN*�����"���L��jT��,�{��Ft}&+2�
'h�0(��F|�?����7�����)Sl��f|����]k��qzUP���������~}�����t\�蘏�R�D�+��l[΄"^x�
�0&�ه�MNt�^=?	��{��Ҿ�6}{&����;�J{.vŮ��Խ�}�N��A6d9׉`������B��y�t����FͿ�F� ����P�d����=>���,���+l~�)mu[�"r0H�������m�pX\J=)��m~
��:�=��5��y�K_�.��<��6z�p����2���b�i��l���
<�CGc�PK�m���sb�Z#�>㟸��"�� �yvo��{Yŕ�\
�m�<��;|���H!�����*�ε�<�{��
~,K(Kr_k�/[�qH��Wj������#��'�S���؏���"�2:��7!��u��~F+2��v6Z���`��,F�/l�o���l�Ԇt`Ҷ��i,�K��jJ�E^{Q]R�kn/��},!���n4�Wz&�]��?(�^�l�S�J<E��D#���S�r=!�j�ٍ�l����<�z|�<��V��l���� ��Okt9!{���0�	� ��\���c���l
5 �L� �u8��8[���ÝG�N�������*��_�X<��*����g�ʵ�cɚ[�X�!���#��iS^�̸F_�����{\���~��+Y};�gv��Fnxx��M���t���XlxV64EB    fa00     5c0�I�����4F�:���9�,�=�M�������-�����T:I�ՙ����	[��~%��#�7}�Y�?�^϶gm;��{�@�Cv�xx�o����r��|�<('W�Q��"S���u��٢R�?A�풊o�Q2�k*>�[�<��I����|���3��	�4��.�Q�V�up�fͳ\n�7��1�V�n�+�9��˼^<~���Z�%uGd���)�A�
'5_��v�Ɍ�lȵ �af����0�*HN�����g�9Q�&W���P�W�h�n^W4��>��&�P9Vo)��7P1j;k�8��f���u�Ӛ=��e���W�[�eIA�S�T�ž}�fu���W�9R�k�c#m�
&DE��ÊO.Q^�'��� |�w� RS"H˙�Sa&0�hŎN��H�ȹj4��L=}!IWmэNw��p[ 3D����?����m��� �w���i�Н�&2���Uj������la��2*�љtp��v��G;N ��VӋ��p���c `��䶁W�&�v��p	>#�L{�G��"��(������ ��i���Ꝑ�}�"�0L�{_	�U�g�q,��/��[��I�u�B��R�̚+��n�3��E#�*3#�E�Ep'���~� �Z�ΙE��^����I��T���NV�W��bW��_n�*��h����ڼ��T�s�6j4!A ��)�h^�e�ץ��w�a�'��ܕ���B�1t;�Α��ꑚ��Q×z�+�|K0豔,ǎ�(�-�S��%9�u��2�)�p�W�3w���ɍ8s��������qO5��儮����C�w�يe>T��1=�� ˚��/7�
�3^ �:T��&�܂�RE��0�l�������#�gkTY��U��@cN���O>&t}T����q`~yl�ˆ�"��.�c����"���Cm>L��aT����b�W���/|*����JT]G��Ө#�04Z/�s�*�^r��:�fnG��S�L�I7�Rm��oE��uX_0�����&ءSN�n$�
�ϳ?����N��Z�����/�)X.Ӏ�p���& �>���u]�3�u�P�^����שzU�7�:lz�_߇�.�N�B�����ӹ���IMy����خ4���̥�{Z�c�Ǹa�XZ7�[S����\}�-�ʧS="Sw��z�2ә茀b����'� �y��[ɴ��TD��r�vJ^1��]t�T����q���c�(�#�8���F	|v'��O�j���2Q-�F� ����x��Yl������Dp��K4d�$K������0����<�Sv�0��D�n�70h�=^+O��7�̰� �䷴��@#�7id,ێJ�ʆb���!Z����d(��f���T(����Uh#ͮ���hB4�Z�@�T۪A-w�
D�����ڤ����.'�>LgSXlxV64EB    d869     bf0���y���aS�����@/�uPo�`&�$����a��K��o?k��I���v����3.|��B;�+�I)�j8�F�i�B���.��)y[ѻR<���l0���������a�`h���}c-�������r�~���꟫��(G�R�6�	9�yK��iGG�2�����W�S��f�$oVk���i0�����V?i��_�6B0;�%/X5�����2N!�0c��k�!C�	������Uԡ�N���t�ﰭ���8�jaK�Y��b|���C �W�0��"A�L�T
^KȨH���>��|y�vBrBǕܗ%����5Ȫ�<H&A�������m���������z�-�*��<�*���Dy��@z��u]]��NˇN�CoYK�
�^.]�/�VX�'>�P��$[sw�12����||��������+`�K��x>-���k�T��@!��e	I[�Kk��d�2���ljⶔ�j�O�
wܰ@��m2�?�P�P&�\w�Q� ���	��CB��������#�]T	�F�8�k�.��Rʆ���3�1C�@y�:>,�t2�2\�v.�*��t���@EX,h�8);��g�q9�".쁰,������̨R~�d+r5n�z�ҠG���	�2�ߓ=/�����T��r�����t�cM�.ɭ_hٛ�?��t�wu	��c���o��^�ƞ��pLht)t��+�M�d�*��YZ�B���n/�)���kH?�_�}��Z��]E���p^��d����:3��{ɤ�4�֓�s�@��t�������/����5����vp��}�;(�&�1ye�t�ݦ��_���4*D�9� �J��\}��#Y�<��D۲�z��-}/���
�C�&��)@;r2fJ�B�C��CY{�����9hЭ���XZ��&n22���FnJ����d����R)u�A��Λ�v~��͓��S�����e��@��Is�k�
���+�ߌx@�2�CϾTh�.@���h��8pg��S�5��B�F�,�
�7��k��o�hk�)%��/kM�]u)Ŭ~y���Q��� ?��G�w祴yB�Q��
M¤@AC
�L�J�!�����ePR D���H�ھ�k��n1O�Ӣ�Y�.��6��p�X�t+�Ӑ h�㣑4�����>�*�G���~��Ǉ���$�q]2.��'��Ū���K~�Sj�{'}\��1ǳ��e��KU�?vM�'T:�u�	H8��3�a���� ������A��*�	�x�"6��-��Ƶq�|�,��<9�$�����r��&н��@ͼ���F��������u���娕,�/�-��4����E�+�_��tg�J�~h
���B_��ZOآ�6���Z׹nrM�j?�c+��Mŷ�F{��q�dT��0\D�#ŰzO\+bUFs1���O�QmAG�t2g���l�eػ�[]q���.����'���=�C-�3Z�wzGX���!�='ۯ,�1S�J;it;?u+���g����\1�]˟� &�a��6K�p�F��?���	ژ�ϲBӦ
H�\��H��Ԧ��zX�\wP����[M���Q�xf�|��q���xc��j������l����T�c6v�bƽ�	��0�i|P�3?qS��G~~7��zWX߸l�������G3�Z���hH�nz���A�i8�P=j1Elo:9×w�tB�4Zqp�dؙ�G8G��Rx�g�d��4*�H�^����IHQ�����,X�;�j����m�-���zjvj!��㯙ZhV	�^<>Q��\����ВK�1j#��_����^Z���O�)ۂx�>���x���4�Ԛ�l�R�����	���?u��Mu����i�l��}ֿ�%�2�3lY���=�G����xu�
_���|�8w�@�_ŹUe���1��W��ޱ�,�i ��5�y������0�(���6F�`�#�"s��+����^�r�j��I�I��F#p`�!�5t�6�@���(���:��X`؊z.l!�uf�RY�@�"(��?P��:�]}&)�[	ax�da�L�0�H��!C��|�Z ���˘�S�m�����r8:&q���d����E�g�Їԡ��K� ;t��A[6��>_�T�"K5�n̥�z|�[�9�.�\�q���>m$�+���/�;��V�e~"�6HV�V�'bK���K��U�*����#�C���4���O�N'��V������{�o�X�����+�c!.j�8�jU!$X8/����/�L��;j_�Y��O��#
T�c��+߰\B�|���7�|�%��蔶.�&ܧ]j?���E�8U)�s��^�x�}C��-z.y���
C� 8�L��1���m���oC���W�w;nP�D[���)!{����.ޢ5��k!ݔ�h�J�'7�04 =�:���?,>pG���Ie�����q�^;�=��)�%?�y��b�[��.5X4��bh^��d����6K7p`�{d%'/)���F��N��)O/_��K��U�?mL��0��@2�`J�$=z
F�,CD�v;8{a�m燞}ob�@�q�@�a��bi=�ߗ'=����z�W(=�ΕO<��dx/���j%<A$�״X�п$1�4n/�ӻZ�xS�ϲ����Ӡry�s����,7#O[���>=3� 1�!e��7%>R������H{�*2�3 �)ƛ������#��B -�ݓZt�*.->�kq�;�k��	�_�_.����g��P6���^.�oKB1�2.U���$#ѪH��p����$d��.��v]j��QpBS�{�iD���+���D�9���z��9�K&e��/w�5*��R �=�?/I�O���B�m�0.W�N�Q饴9.6m���{�Ĉr��&oV��U��0��������*)q�X?�	�P���\k�[��q<\�3"��