XlxV64EB    4876    1100�@���ܴd�~�S��0YqI�r&�Aw��2 W�%���doǝMS��%UĿ���}�L���\1��Z
�i�5Ѡ_��T]@��b��mz2ͺ�i�!w��s��K kW-����C�\c% ��n�R�[(�:ąȘag��r6�������o������,��8ꎬ7�����!�~6���9O٧.�L%���-6��ɸc	�����q��Q��P���n�o������> kiY�&��PH�.ck�P��^��]|����������{��>��L����}	o(�*�	��7z'����7������qT���Y�:4�L��Mݵ+�.{&a��M׿�:��>
Fp�*��$�pr��
$���홸�Rr����t"��R�%�,�_�)����UP���	���L�S�R���#G~^c/�:WM����4�@;$%�*BCKO{�� ֠��t���l�_�M蚣9J�
Ə]�c1T��ӹ���ŷc	�u>Y��t!�m�L��V/�o��(Z�\���~9K$Ro���#Ow
~�w�,���1v�Ld�r�?��4�R]�I.��%o9a.K59o��5�{��:�|�`&�k(�(io5��f��`h��S/��2�y�������Q�)&�8T'�-	�P�˹t�wI��'w�$G�"�K� 22�s� �w��}��=h���d����v��]��E�!eJx����v��ĲȽ �d�S�oA�Z4kz��Q.[$o֦���n�~ʫ3�UkX&g�W:tN�Q}Ҳ��ԧ�VGY��3	T�%9��/(�:9�j�,�B�G'�e��W�B�h��
��:�W��V�n�&r��ơ��u�A�'��8v�g���M�0G1�����mM2f������X�`Z`�^���7�[b��цN��լ�l����>Z���h�/�(g�Ș⋔�����A�J��i��|$-9�c���Fe( ����+쌇-�9!`��,CD
߶�����	2}���4t�!�O^EF)�
�|��z����N�����Cp��_����֨�E�3.������hT�e�n�	0�wg:w��9CRz��-�����	��t#�â����ňx��~��u#D1|�Ui71nc(�1��~��V��I�j�q�!��]�[/��Pd|�G�z��nPyՑ�r4B����"	ɢ�?�|J�hnJ�@�o��	�%��V�˷̫�`9��x���H�p�/�nJP̰���$r�YX�`�NǤF�M�L���w���ø-v̗�|�4��@{�$� �C=~Y:�0��ɵ����t��K�f���Z����0�ۘ�q�+}���O��)��������H�LN���h')�"4�Z���7�R��R�����i�/@ǆ�T&O� �E\�%LIIK���Mh�JA8)d��5����}���b�k�� >�IF��T�������O�n��Lˆ�g`j50�ʚo+_��:"��F��#���~_4b�� o'�|C�=�]Ϙ��-���$Ä^�ȫ� �2�
�clO��6B�q�-3P�%�89�;��_FB��C����@JI��g����3�2���ܝ�'R-�4Çe�,��߼D�3ܐ��K��ܶ�%h�����)-_� �K�m�F�E���j�Ǎ�Yu��>j���kxn5����ǧ�������iS���L 4`_�@����7�k}��W�S.�`�wƠ"��A���|��דQ��{�K��t{rkT`̏���c���-�c�8�蚚t��- �����s��+�I�����qV!���3���>T�?���$���D�sWt�Q"u�':Y������7B?�@8�A�i��XچU�#��Ӡt~�A�Wp�������T+��&�ݙ��ի�A?���0��(�7���jh� ��ݑ�D`,�	�9�	�<��5;z��
�d{	���)3��Eϙw�e ��������L&����%��˺T�U� z�1%��G]
v:?��ݭ�8:� �L�(G=qt\�w�y0Ӝ�ў
�Aݲ׏�O�7P�#����L��eG�E%�X�$�j;?��3`-Yݣ�@� �7��"�~m%��"����	�&!����S|X�K��#�l����
���f�XP(w�gl�	�m��������\����v��l�+�����G�O�8 �9AfP@t�{̱9H����ף"��,��?��5'(�E�E�rx�S:�\X��'z�?ی$l��k�Ρ-��������WH>"�4@ �D�ա�3�j}>��K>��F�beu���噧p��Mh��V֘�t��[��u%�ݼ��IFF'��X�2�dTF̫N��*��6Z��{q�I� ҳ�4&�.b�����cz��/��$Į	F�ѻ�8�,p��������^��+���e�H�qІh٠O}K]��ĉ�����)5��t�c�����毠7�7y����k�{:�T�<��45�y���%乞��,==��XΒ�*�� �B�,H$�Fx��@�q���3�j֌�H	ݥ�X'}�ʒ�*�o���܆t�T���Y#e��{Cg_�j�NT�7���c��0���*��z�^����:UY��wc)����Lt"�5Q�Rz�)��&~
��H�B�w%��ẘ����_u�8�f��8B���-	X/.��C��l�)��Z�T�z_M*��B�6�63R듵�#��9}l�a{%������,��hm[Zch�UA"��:oS�(��n(Hs��6�I1���I���o%��/-*��-Ww?ވDSQ�����%�	UR���;hm�Î�1-�_�/)�7ʺS���J�f��SC	���Q��g��T��B����@�P��g�(�w!���S��ڕ�0�Ӹѵ�e� e����_���Rl�	��5aѹ~(UY> cämp	��M͏�|���4��M��4�wa�O���Z�EƛI�!�`=�yH��b�OU�����:剏��a=:"�.�
��n��A��W�5��
A��'��\C�Q�{����љt�4�S�wu�:�\>w���W,��e1�':W��/�<+��#��p/�{J����b�2~p�����dl����̵�[۰�V�Z�(�������~)8N���o��4&�|��Y�
Y���U�D�i�ZP@�^&���	������ի(:����?e��E��$���m{��9��b]��Jƪ��n�͂Ey?���?�?�m�֭*��4�,�ሑ>�=2ƀ(�u��p�O��;�[0�I�Z戮����Y:��g+�5�D��Ă�O��w�����!�١��.�����Z�_�����d{�^��+
X�!�v۩jx�/F�g��r̋W
J�c���!�#Tlhi
HM���$z���?�`	kٛ���i�>D+h���~a�ɣ;�[�ǘ�(�����*��pL�9c��'J��ƒ��Nb�9��S^w�xH�g.�w�F�l�n
܏c�.1-�����|�5��e8[�5��X5��&�I9b:�_[c�Y�5�W�l���q�n@�H�F��TXjs��Ke7_mw��W�.@�6>�3��L�ӥ"R�p�D�X��8�EP�F���zQ��t��2�lc �g�:E���:5RD8KlJ�g�	����|N�_]�9;j�mu�F�:3���>�X��r.�a�AgQ'Q�of�::x�=�:!�_\B	{#���l/B�q�9h���$�?���+��P��)�^]�:U��#!Ū���6X+c!���e�-��@���U'���>�+��i.��g{bThO�@�	ʀ��C��*o��&wAs,'�o�`"���}�`��ZuG���p�4[��i��	qt����A5ZbP��U5���6H��1�YM�%붯�I�k��:�9�˚Sgv�d��t�5!S1N�V!G�n�N$~�B��_�@�vY�չfR����yK��H��Q�7[�R����	oq0��Y� $α���_�"������:�6�+���Q�D���[������Q0����4�/0���c�,`�η�<����'�v��Bh=�ץ����W�eW\����1���Σh��_�"W��>j�VN�i�~6�$Ͷ�znh09�N�sI��v�D��Σ��.�̟L�o��Ơ���������B��s�7�� �$��i��0�� �ׯ��L��0)� YJ���꽁ʹ�����Jbj�xf��B/���Ac��4���X �q��3�Y�N���!e���