XlxV64EB    4f6c    1110r�߇\cD<�v��^9�1��k.y���9��;X�vd��� �δ�e�?했~�^����/ �Te ���3�d>�>������'l>D��<�����b��v"�����`*Զ߻+��ک1t�ǣ$��n�[NL�Q�ձH/�̜} �Β��{�	�"MBn��`$r�r��$�!���t��+h�uPG+T���-j��F���g��*<:�g�F<d% �k��׸"��Q	Y�͖�4��'��#���AhN�1OC�[�6�\��.j=bê�
񉧅ɖ�b[L�����@�#}�x�o:��վA�_����gS������ؘ8њ�������L���~�=��A���a�Dû��ѩ��p�fʋ�)ڗG�f�+a����G�亲��h"�m+�s�D�0�:��.��ۓ!|��'�u)X�4_Ǻ� �){�^xt~�RN�(�8���7��㦔E�K��ی�&��2bh�M�d�q�`�G�p��b�`��+�?��qU�W��s��B�M�|]4��5#����B�،�=��%%r���kx^�g���33���'E�`Ӫa������H��O�%�z�S�FF��+�u �y���K\��+��L�cP+����6PM���Kw����1�Y9�諃1�����F��[��S�n�.٠�����:�@w���3i����e�ΚLJ�JJo2�}�k���5z����4vx�
���N��0�7�k�C�?��2��B�(�
�Oܚ��y�\���r���\C��G����O���s�.8�p%A���҇T�`���Ӱ�3��L������tӛ��H��|B%���x:TTF����s������0)\�}�٠	����6`�+���\�L�6��t�%K�$w�Bifn%)#�L��=��	��W�A��]�Jt>���+�䶯L��P:����;��VFN�_-`�C��֒>蠻ھ��bo6Ѵ�_]%G~!�#;�	&�s��e���Ŕ!9�-�M�O^x��8T�}�����)�R}4o;vg�+��hԼL������%�1���@p���px��TJH����0Pr���
̈��H��zP�n$�� ���y��*�q ��O i�Y"����pO�l2��V�!���<5���m-�Qs����F��؏{��M�/_�(m���8�8$+���k�Zz�%m�qa�"~ \-�zBN�>��	b�q�q�(���c�?�K� ?��#��F=E���tjo	������m�q��>Ǧ� �8��;čMZIZ�^�&ur��i)�%�i���r�x�@����'*����^nux�����"[�S�]?�9t>���,�V��33�ڜ�h�Y�ef��e>Ì�$��2�����%�R�!�dV��%ӻ�
H��*�'ٖ��*U�=4b��[�����C=��C��U�����J���v�e�O	�1g%U��viʲa�t��B���m�C~��#�𾊳��h
3���KH�=->j��M�C����=����bs0[�ID�B�����9}w/γ�f�PCW����CZ��E�M��-}���ks�ˮV���L>���c�g�k1.�"�� ����c��*��]�D�
0�Y�`�9 ����;]�+����<�%D�H����M�gב����_���__aiB����v�(����C~i_&>W�W�f�Ĥ����,�Hc� ����r�����	%�������,���=[o@,� ���j�ݓL)(��R�?Q ��u�Ϩu�X��=�\|W?�+�!���F�z�ժ��l��� U���m!U��jfOַz��璿Q���G�nJE��^� H�6��h�{�ހ���F�i��L�s!;x�Ȓ����K?�e�E6.mK����2j]����U����ƖP��`��0Yc�#�SyM�)�4I=�t�=wo7_�%�
;���=�U��P ��=!���ֵAy�o'9���xu�����k�?��el�I#��G
$�̤�5���rs3��<�wjV��r7ë�bV���~�o���U\9w��e�ͱ҃d<&~NQ\�B���j���?��)�F#�&D|��QR����װ*zރR�=���ҿ��*�0�R2�@���sƧ�pj>m����Q�.�fH�MI��"0�ν��>�uq�p]�/#���Y�ݞW+�N��(��8wc�g"�^�Wͻ���B��Z;1R� ��g��P��),%}�ݳ�.�����2ݼ����-�'��XF�D�*f�I͋8H����˯6�n8�ߐ��M�$���+Ig~w:p'�P~�6��_̷Ѱ�V*��\������'n���ƕ��� �cb�:�d`I>O;�P�{ɟûԖ�"��u�]?0�5ů>����b),�%Gh˂�)�����5����A�}˟gՒ��et���|t��h^��y�AA�}��{�x2���ƾ@�#�f������5�[�ђ؛�V�{��
Ӌ�M����C.�1 AZl��Ñ�N�*Βhnp/p	S�Ww�aw9����Ř�?�
�W�7���%M�m|5�F��ً�!�*�,6CZNL.H������j��y���,IX׮i�R�с8�%�B�4�<qi��	p=Z����R��i}H�J�=�UA,�f�PB�4��c?�<����ƹ���F�M:kF3V+���S�G7@T���j��W�NS$N91�<�X�<{�4�u�fqT�B��o&"�gY�NkS��!v�ŏV�u�0�0��/�����p5�w��6�,�r�=>�t�L�uA�(yQ5BRW��R��X�`:h�D�2�q���n?�2�N��p��W�螣>,׳dHq���Mr%v�X�뭏�
M��a�/}Fa��ը5ޚ��=�g%��K�c'=�-P�\�����d��U/�`̏�C	Y��-k��o�+���TvȅQB~��
B0��2j�\-�T9�Ϙ~UF|��,�L9lǟ��y������MNQ�Ϳ�0�2m�K�oƇHO���[z�?���=�)?1��fVP�S;qA�c:��0���K�4n��J(��>Lg�ڄ�ʅ��x�c�\:����5�J�'�p}$����%�M�"��*ŮI�A}b��?��>c���3�\7�������ι��E�]o�T�k]��Z���k��*$�!��Pa�i�>�J�Ȕp�d��A!M<�\|^��q���0�ne�%����~p�s\XӬ�X��	rZ���a���Y��G���(骍�y5f���q#��[�2�$�ÍM�0ٍk�I�>=G�~<?��k��mvm�Fy�"����Uu��*�'"��9h<�Ģ�*�z1�MdLHc����Z��g $ 	���貨��$�M�� '�(_��#��j��l`�e�(�ǆ���D�̷�0$�Z�;YK����9���p���RUŚ#���,��.8Yl�:=I�e�{�k�� �������u�M)+�z�Wy�}����,o""/�vi%��8�W.셭M/C��m`����;�>_.F�G2�I(X^�8��k-�R�;w@��) �9�^�GQ�5b<B��xJ��2��{���Xch�ᤃ�A���lkB�n�(��;$��!���Ppaݏ�v�'ðeYT��%�Z�e+�Gc����J[���I��Al�?
t/�r�m��� �i�ݓ�4L���̘\K>�x}��1Ȭ�'�p9�⚛@��I�g�ᒝx��2dN�ps䙉����P�+3�9��mۓ�]�]>�kDg �X�3��\2z���"�)Y�du��� �YP�8��Ԕؕ2��E�����򖧊�$��)��b�8C!�ؔ嗒K���3+W��*=�+n՟�Ѫ�%В`�Ε��d�/�e>�R�8��}j&�w����Q�� SI	򖣎�2��󎉠�>�(�,i.`JsQ�up*xŚkW�sf�26��M{��P�O����%B���U��(������b�Bo��NE&��9�K�yX2)�O�-�1KB�����)|BO������N��F7"W�#B��8OGEbo�w7���?�$(��ot{��{뢷���U��;L�è�̭���G5��in���ahC�	h ����/��Fa�����_��!eﰨ
����oIri����6SZ���*�)�q7�I���{�~]}������Rʡސ
��S�ؓ�%��> i�����㐵'*�W��מ*��D��cް�uxB�vD�>u���+�#"c�r�mܫ#\�ds��@�FT!��zՈK�w�D���&.��hZ}d|<j 