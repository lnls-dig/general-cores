XlxV64EB    3adc     f10P(鰉�˵ <���rlK�ܝ33���5�#�뎓6��W��ƙ����e�JiZ"���d�A�cn؟�>���cf���%x�UC?I_��O����.�1�V@2:a�����H��)�r.Ci9��m�U�fz%�9?���qzP�f]#9� �4=�����#>5I[+ޝ��2���O��.J����AY~��%c�ג��d���h�GOkW�i�O��|�(�h�,[D�������0�rm��<~��vB��ɝd�����̿�W��X}̎����|3����a�C�����W�\rv��_b�_��B�:=-I���PǌވXY�]���?�l����(�aA>ELB���A9���`�>{d�7�*�-��=���� �۱�\��2j��X�H�Z*��R���D?I0u��iG��"6��:5�ƥ���ɀ��E(!���]cS�/��K�.)υeg�5�&<�q7�B�]x��[`�_��*�J���)bDj�lrEnE���@�8׀YT�à��sC����O�4��`�)̦��Ϫ�)���"FH����t�	c��aA���^F�����*	L���p��nO�jZY��|���#���^割t���<~@܎�A��ވE��a;��oƺ9��[`���vn�ĝ��A����h����xT��r�~8V}ͳf¬�%�#���V_��Jgi��}�We���j}A?�=�6G�c=�X���h&VI�
2��ɦ�����nJ���e��O��&c�lB9���Y�yv,�a3��;�!��FX�%�|5��z/��>C��|�lʬ�G����I���R�Z��T{�:��?͸_ڏ'eLz��Igf�&�/2	�@��O��ǽ6dD����M-�L�N9LF3>߷=`�Y蔐�ۻ4�˽�p(q:�I!�H�>���@�)JAW	�aO���[� ��~5��XN�I�%o��r�嫉�qX�s�~�_��M��BΕ2���ᘿ~4�C�+�&�zI��`�IN�/h��>Ȃ��%��k1����p(�(��D	H���_�o#�V���z�`hq��"�@`6�8s���*�ʚ��x��c��T�y�V+��8�͈:��ɗ����öIұ@ȱ@QD�|x�8~
bDo�J��9�1v���ũ����I��9	V�@��6#L5��w�E �e=>����5��B��7H�*w=��9=�5��#$G�D
�
�����4�./k�m��U�\K#1�'P���a ӥٌa^�ي[��^�aHw��WQ��Y�x���@w��?ġ���qҀ5���VA2��g��磏��D��qQ���\[T��3�n0�8�(W+[æ��̵�\�{�~����r..�z|"�A� �`�e�Vot	���}㰫����n��g�g������ڑ�[�����*�#��>!S�!m�b�^�ykt*�l�1쀄����<b�d���+`����㹠�r�����d����%[B/�	���\���.L��d;$����I�*]������C�,�^�U`�A%[�=�۶]m86n�
����0����CL�q�=- �H#l�:�q�%��\�ΰJ{�m�����C�p����0�X�&�"s�U?X�m��Oc;{���:�"��%��i��cז�}����U(��eVb^��+`�1^LH�a`�m0�^~�닷D>}_q*/�w���y�O��+�-\,r漹Qф|A�x���}��>� 1��%J��s����J����`�X*��*������=᢭?���Mw�&}Er2�6@���dƟ�_�:�O0[Q�/�iy��w�*���l����Y�JH��N~��]��D����c?�<�@l ��*~|x�:�.Jɒ��53dxe�bZKq�~�h��]8��C��K�))͢�/x���p��-A<�(⍀���^M�qP:�{��l�Q��!Wv6�w�p��B���v4��e��7��;h���xrr��\�;�s���i��+.@*�36��G^~9��ưrqvyX|�S���	* z��a|x���B��0��� �����)-����_�-S�v��oc����x����qá��؃p����	�XVO�J���I�B����E��;�����`-�E�1k@�tp�G�Uz���׆ou+,%׽po�;��k�
#���������a�$)�%���*���7Ч��ejF7 aB�-�M�e!?��@�����A��[�TѤ���N��s$�@���hD/��ǀ�_�ޒ>�ql��5ϙ�ϱ���$�t��KN��*�4���(�ϪS�,?d�G&I���X\�^�H����Ö�?U�đj�>�z)g�e;`��=���n�^��ޮE���^Q�ds��u؝I�RE���{�~�(r1��y�����VQUƣ��p��.���7ͅ�^��-�ÿ�M�EN��*�Ê0��T+�\�w���c�6 ��J��B9`-$q��7)���
��s{��HA��1�����qE7&|-���z��A��ih�]?���G��f�HqL���ˇ�I�Ļ?pt9V����
�y�n�N��x��\�c��x8�0�*ڊ��_�p�;p�%�
�ۍ!P8;�Ms�2�5���1r#�W�/f&aP�_�k�>�
�Q��"�Y�B�]S��ʸ�_��/x�5.�!��j9��L��,w]�T�\̠�Ľ	(1;/�FR�.����o��nsy����֎�e������߉ �>���N2�!!ǥ^�Nɣ0w�-\'efWx΂|a��d�l�6����UB���9r����ZZjԐ�3�<S��_�"E%�4�ʎ�9��XC�g�v7֨���%\��|��u�w��!�T�j��^:��+%&�!'�`͋养��,��u��o� I�H�V��9G����M6���qa��a	�Sw��f)#�#�`3>�@�L��8ߠ��v=����b��t�7u��y�|��TM��,���{��`?�ӓ�(�E#ﵛ�_�>�K8`�M�K��U(ߞ�2X�dx���t<6�,D�=BRg|�V�5�{��o����Ս���S��$j��ԧ�zW5�B���G�������g���Aƺ\��Q`�7��	Yw�7�)���c�s6��p�
F0
��y~�՘V�,x3NfO�?3����;'���^])=v� B��M����$��r�yXmᲑ��O����A�jm��M��2n�����9d�Ў5��K��}�>�K�'Q�ܳX�KҌ��Îa���y=�
J�p;�[�h����!��n���ۇEuvd�=�������������ix���<������ Y�`]>�?쇡�!�%���`{s��t��luJ��%9�^�[�i�?n���d>�ϋ�����毋S�+�\��2w�I��Cph��лJ���\��<ھ�8k���;&��l~�3's�*��>�,�RMp�UB���N��V�L��Q1��jʀڹ'�q�Y�<�i���ġ����9�qB�P5�%���`�&���)���D*�D"��!X_�ꏲ��Xmrc��&��/�b�5b�y��
ڭht�z7;գ�����鎹�uj0$V�B�fA\�iY����%m���}K�}�ޱp�Ö��u|�&�G5��M�?���o7TX}N�T&lL��s)��i
����������(ɋ��j��I@	��
�iH�--a�Ǩ/�+�0:���C�R�����\;0���E��Hk������pł�9�oE"�<B�Ԕ$���/�h���Y8�'��UP�>�C&�8��@�ea���P:��&