XlxV64EB    388f     da0?��a��b��~�1�+"dT_zK�vn�A�jU]x�:�hz��S�&]�gN��)mL"��`��Y��2[��5�H�[v��m[�~��^�����:��C�jEF���]��gp�*���ȸA�P)M"�U�s��a0���/��4�����;����iz���!���(K5Y�ަK/��������|��R���_�[x�7WW���������>�����
������/У��w�!��H�(Jb'�<�*�Y�O,�'�R�MX��Fs�`�����8���b>�@���R#���(%�P�om!-x����B+�jn����_�X��s���ު>�y%\���" #=Ahz0�� ��n'���4��6W�u�>�����I؄�`'M���?~�Y�=�w>������s�ҹn�2X����sB&kN)��8���	PPQla���B�d$'��:��K���
*�!��9�Z;t��
��a��x}�9,W�z�o��q��P���WBFL8�q�t�P�\p�G�Z߹�����@#���Zo���If�s�'�a�޳Oc�ED�2��L%+']����!����[�b��i>t#�z8�5հPWW?�����'�B$Zj��8�P^�V����(��a# 9�5=At��a�Y|��#1��o�yx~R�R��J�z<����؆E�����|W�����'����c0�j��g�\�%'p|'�Ɉ#���f�6	��`Dӂ*���nk�G<�"� I�_�Z)��|>�.*`�U宻^�klwPcձ.���D��l��5�kE���h�:l+=@�P$�g�v��縓p�j@��P ����Bq����mq�u{C����3+^��l�~S<g���L��GA �J�I�/�0o��O|냩���R�6�p��A�j��O�H�hw�m{�Po�����d`9��Z��)��	�7Mc�tSi�\�+���� ��?O�Mn|>l�0��^z�ҁW����{iE-�%���� ��� <�pФ��I�2��;k�>k�����Bm+᪑�T��ܯ�nD�ф�%N���dO3&��R���-Cv��F �U���H�Zj�8�T���cF��U�bx��uo-��|������t�a��o���YY�·�F�$�%����&�U���>yP�*���~�"hN�{�5�����ܳ7����t�$e��s������
�_0L��N�88�����+6�G�Cp�R�'����K�}�|.���o*��Uk�<b���:��i`z�������b�{W��>�K��6�ԯ��D�]=�y�ėde޿H�á�=9]�"���&��:�cY�C��p��mڛ���S�����A90 �1������X�����b&�:����z W�)���t�JǨ�%;�GľN.�J �h߷��Nf�T;���#�S��H���%O�B���/���)?me8����¼�� �&=�cM���R7�C缡+����H��&�	����s��M���Ȕ���p/sߖ���%
G�!t&ݽ(9�ϧU��m�<mէ�3yPi-\ʇIj*h5�����"��{�YeGm���(\�H��7T�Q��m�� ���iI���cy!�w/1,>��N1�������Z�qi�ׯ0j�q�:�9���"G�HVc=!�4Gɚ��2�K�������1l�����7v�{��Xv����/���+��^�'�<$���D��e�7���>�&>C��M��>�?*bYA������F�*3�Ǽ���,y�hE���+sdT~����K��O6�6�S�93�O8s� ��
��X	d���,͎Yx�L�����k��?�`{:��GBs^����BG�����Տk��Qt��������V�Ԁ�?�@���)�ZJ���ּ�ߓ���=""�̗�z�t��)G��ayx��̹�!�7�*����Nqm�`s��x�a�Θ�H}�Վ�wY��5�|B(�u�H�ӌ.�}�����'�\�"-;������]�K�p���_>M���À_���0+7�XU��ľW�;�M33�>�!�kyc�La��k��t�=��Y�-�B;1�s�z���LQտ�7�U�n޲s�cBxu�q�Z��hE�X	�V�$� V@���<4k�h�k�!���VLؾW�&����uĽ���cV�NDZ&1�XƗq�m�p�ɅF;�iT���Niq�+ړQ�n���ޅ�l��hY-a�N3��R�+V~��n����A�B�0s\0�N��+4(H��Ŵ��@�];&>�����(d�hc�@f��'��`�b?�W_<սO;�z9+�d��Ĥ�_X��޷���^��?8U��)�����)�� v.�'Q���lQ�����,�4.L�'x��J1�ɒ��/�,�� ���8,Sk��ϳ�<����f�U3c�0�m�RU�`�h�ԟ��a[b�Lx���45�n������sƚ�A5��Ο���B*(6�z�ݢ=3k:R��Lj�E�Ң�Ѻ����!|�)�{��M&8v<lH� ])Џ4�m��H6�݇].e���>!�:�L��'�0L�MO������O]OX�X���K����T׍��ЦOB���!ܼ�<O /�8������ 8>�y�[�5=�WU�����z�"����um�* �8�����+FW�~��B�3�'{G֫>S+$r��\������[D��H"d��(��fV�����-m|-���a�x��}��9��
ٻ�1
|.�Ӻ'�t+�]|��\��~�o$!0>b��<*�(n��c�#p��vyle,��\8����X����a���X����E
��l��B�8`�����$�2x�v�5�>=p�ԕ"ˬ�(�gE��;��rC$�b?I�o8��e�l�.�3�TǞ��ǅ�/��P%zi?D��''_�9�Հ?K������p�:�Q�����l�Ya�ZI&ԒY��+�o%�̼2��c]��َt�s	'Co*�7�����AZ�8���_U�v�!�66>ĉ?�K���;ϊ�]��,��|)�U�Pu%�_�"%_<~]��$  ���;�M=X�	;����L�{�y}��)�Adq|u)n_Vξa�O�c����/ut�N �<��Q��1���9�ą���ѫ����*��~
ƌ�W�^��p����b�@�9$���\����r�g��,��ڴY�-l��>P������X#)G�Ӹ������4��ԩ�"��%r�K;��>Siߏ�u��ʡVE��>0r 	� ���QxC��ub>��j�~�5��Ż�N�^4���`5{ӯ�k�0�}�����/\�	?���RH�
~�CiG���Gi��������1~����R�0y �0��X�e9����ܫ���@c��@i�Vnt�W���