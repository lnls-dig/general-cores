XlxV64EB    af5c    1f80Te0߳^��8�y����k��,C�Q����7�e7r��ff勻��Q������3Q6q���r�������Pn��j�"F�X�w@ܢvY;[^]�	ՕC~�5�T d���
�D���Z~Eb��Mc8�r r,�3,��9}�Np:��~���9��u�O�<{�	>�g�u�8hxOd�U�R�^�O��Nx˨o�F�vqH� ��2Xv���
M�j�K}�^{A���Dy[�"*�{���{=k��س{
Q�,"���Iؓ��R�����,e¦��AU�\r��L����sDNɻ�UBU�t-X/6T9���Zȉnyq�G˵��79
H�d�Q�8C�n���պ��7�ʾL)�������m�O���
a=0�R�����y�oDc�6Rdx��M�X�`�j"�(��dR�K��^�C`͈��D���n���h��#��e_��B��`���%y�=��]�{� �}�O����J�����jJ�f�А4I���Y��a��Bp$i�ނig�����Mx V��9���vٵ�E�
,�.jbR�,̚�C%<��O�y�u.�Z��k�ѧn�f�����s�\KL��w]����^M�qٴ.���� ��`k�uƩ:�ws{p�qu�_�P���\��APj�o��j7~��o��"J��:�
�������4m,��V��%7�PCۋ���9sW8����!J ��{݈9��Jˡvf���9��Y���G�g�8ɷ�K\��mNM �gE�N~�I���acG��S�H���)�lC�.��vj����;�c����yxaDop������N�G�Oo�������畲Z�2W1�A<��3���ln��`Pt�������\J��I�\�1|�<'j�Y(��?-���Z)?mYK*n	�'}�yB���f�C|��+Og������hE�W+w��-�IG~Z���Q�����+�u��Ib�㮳6�"���}ـ�0��Q�%�.�i	"��[<���a�(va��Vu�Z�U.n�;E{jHRvv���ݗ8X��☙��d#v����H�h8�M(E1����+/�h��)�Q2jo��Λm��V��K4mɞZ���9��
�s�(��^��̀˴%<�C�y��$��,;��,X�n�m�ZfM�3���$m򪾒dZ�/�^��5�.WpZ�Z����ki>�,v���nUs0ړE���E�x����\���즴t�s���Ѕ���Rx!*��(-~�1,)��t��~�oN�����H"��ڒ�P�Fm1R�ݎDG(�?��6B����D՗~|o��'�bw<.�8C� s)�}�b��4Q��i���[Y[Eӹ(	|�t%�@��J����U�7���~�Y�EaE0G�.p{�J�Ƣ�,�����<1����w�K#s��&�
Ð*t_����� �d�"K��P��u\mt�t	�g�9~MOYRpԬR��QW9Wr�˜$Y���3i��}��6��!
Ȱ�7���BQ��hW�� O�8fMv��+�O���i�5���2mfp��57�7�+�_����o遶����/�?�Z��|����V�u�w~}�hN�O�.$�Y��a�T9�����u¥X޵�*qn��k�xy�
xM#F�tF$�
�z��ɇ)��i�'��ۄ�O�b���'���8��5t��.)�F���!�m������cc�BӀ��(i����}|y�p��	�2��]!�Q�u�1�f?�̼��M�� �ݻ3�|�j��EPrt~Z�C�Tڥ��,�Lt��/\��!�E)�����K3e!��KuԠ[����y��&����p��djf�k/$� 	��'Ll�+wt���c��d�9������Ή̙��a�An��𪧪.b���]%������M�n&���۸j�1SՂ�O$�k��[�r�!�Q�"(�'�g#J�J���������,������	D�e�`*?b1��_�-�bR]�n_)�ĭ�|;�WLV��ӯѸ���N�P��{٩0<Df�a��}¬��������:@�l��&�sv�l�ǥQs�ڌ�����~�Qxk���݆�9b�]�S�9t��t s����P��f��	Ӽ�0ɀ�K>/վ�[����i�cc�3�W������d�^�����bZ�W�Y�]�&�D π���*vU g��sŒ;t��qh�
�41�Q���O<�3��M�f��G�&|n��f���(9l��b��w�|�J�d�<Z�������0<,�-�]+��TkO��#뒫
H����p������Pn�|�j{|�����C�Avb
_�8?E�fSmҽή:5���N�+tTW��Q�U�G)��y��_(���s��U���i*W*��Ail"*mr������ݯ�aJ���-���B3����{�CVp�g��J�ֆ�64o�zP(�����iw�x�k�\��P<�la�#yD6���o�VZa۠#*�	ㅓEO�O�M�u6�(X�|�����Tȸ(Z�f�㴨�0� Ak���{��7�Q��?r�;�ρ� !�˗!
$�c�k�w��6��Y�8�%��z�y�L��J�M��_2"&!=`w���\�Hc�G+���@��D��)�^Xƃ��Ҧ���Q���G]|ͅ�u@U`�ۣ��9�mip1����7Wn	eXB�j�c¨w����C6M���������D���@�3U�@�0�t|��coH0#��C�rgʻg��0�ϗ&u����
YD���?�(X��𩖷Sy�!���v�2�~�h���(�;�lS�V�`;�e�^����ꎙ��?�3�a �� l����A">CJ����AE+��n��>�ǤC��<J�y�`K�������d�7� ��,l��n�+'5���G*ҥ2r|���Oa�h&�RTX��-���չ��k1�Ў�a���
��9���a��}L�,�\�;Y2��Ƿ=f��
��!V1����]�v�@�`��.��͝�砶
W�EJ,���K:�66�N��~���}�Aސ���ߡ�1�7��;�?D�n)�m{���l��lo��2Ƃ�Z�����lN 4���t��ݞu_"���1�zp,6�G�;���EP?�}`����~:�#WeR�x�������*v׷�s+l=~Ӂ���>��F��=�R�,n����3��e�tEALdם��=D�&FW���BJIK��ߩL��RGR�8��0ڷkiƺ[Xt�����F�k�_+�g�����t��h{��xU��LhlLO�D<�)hHɏ�~!38�ˤK$�\'��a�6���9�,�A�z�����"�%�<9p{K*�����X��y�ækO��K�_p�$H5�?oUm�h࿛b#�ܘf���+��~zv����8���5�z�M��0���b-�,�'0O������7�6)��z\�K��\�-KEV��4�C�'�b��r;���r
`\&�&n=V��Y�>ɼ���� Bp�axY�]��bT؂lK�k�CL1.DB��h����/7(>�R�����g���S��B�I�q��,AjQ���8��(u��ES4�P[�����c1�4�_��j�Y�&�,����{�+e3�����f"���?�k@� ��Kk��,����7ǀ�z(/c)҄�s ���"�����XF;^�d
����F`���z}$B<A���C~ET{{���^"��2y�p�n\Ye̩L��W^F�.�W�lS+%�
YX�d��ru�ڜ�$OK(fp��E�����E��=З�;|1��8f��1�X�!u1�@�Df�6{��1ۼ!�*���e���hՂ�h����P"��xT+�t�qŇ�����Rԥb� 1>�[����j��T�Z@5�|D�G昧Y'-J&<�@�N���p34MW*�B�	XaI�г�	��oWFE�B0<3 ,\/���o� <��ޕ��j�/x�Xa�p9"!�*��,	'y�w�i�� rB�S�뢏T��e��^�~Y�.}��s��:����cLt'�����+�j������-9�L��d��k�
X���$��z��ADA�K	���Ga�q�'5��ja��@���*�jA8�b�h��UK�Dk��2
n����|�@̣��50���0�9��2�}�慦�8=�/ѭh鈎�T�9M]�*��Q Y���2U��
�����h���O�����P�h�/ă�	٥��
'9Z2�(�����!��47ڭ�r��;�xX�����w]�C�.���1BG�#�l����۳�z����x`�"K��h��Q�oгk�6�]�_�/Wn��Af���N�U�|����BŊX�Y�Wku�[�q�l)<X�E��m��@�qi5��]�c��x�
5��19�-�P�������~{��S���Y� �Yy"�Fh�Q���ł��1����ڤ��H���B�~onE���ښp����A��ѠE�/E�O����l>��#Z5�;�`Q�u��V����O�.�ś"UT/_��mz�+l{�G쳨NԫN���C E�����$ݴ�EKc���`B#�#�4IԒΥ� �����x�ϕԵz�s\`K��0�ܳn�:�.,�D��β�d���"u�w��MF8�.ک�Lدh�B�TC#��Q/q�ޣ�v!o��SR��b�fPI��NOt��h W�[1�M�U�"�+�i_G��l�����:���{�4uaO@�Ř�1�d�B��f��r&��ǩ�$2�j�R#���m�l��;!���x��
S"3����|�C�+��T麯�%˶�Et
���Dh��*ܨo`���ܒ���+F�܌V'S u��Q�'O8!��P�Fo�Oҍ�j�.Cr��MR�7�֧������RIX�LV�b5vm�n��(ݪ1_a$B7�����J�د��w�}�?�$&�I�+�F��΃�X���ӵ�`�襅�$B�M�^����)4@ ���-��٪"İ�7ŦپW���ŬS;Q�r��1
"~~���7h�����6�[�5��d�j��2re�M�dՉO~㗎��q!�̩��4���k��=$u`�[���-ϝI<��}�pI�g���{�ɺ_1 y�n��r2�)�4�6O���&XN�.��h�9,˔_,;z&�l	Z��A�ŮA  r����.���n�������4��� �Q��c������)�(>�CGN@ы^�Y%��u+"�nO0ۀ�������C��>��9�ނ���ze�G�l\3c�L�g�M��jn�$t;b�(����a���glo4�t�/* ���� 9__��L��������������9=5H��(aL��dn,��)�=�[*��7����.�Cz����VYg5�#�z�.�o/��So4����� � ��WuJa�ÞFXs!M�`�l�����V���D�����R5{��g�RqZ9�c�8�sy���J���%�ݰD�B��?�f�5y�y
C���=+�D��)/.�-S�𗡠�?�ڷi)v�&��t�SN*X�f�N��"���<�1H�:�Du�QjW4i �x����B8�#ޝ���9^(<��ET��3�G�>>�L���:TV�6[�τ�/��WBҠy%�ߔ�\�K䇿Z�*p����ww5��P�:����q=�-��m�nj���)Am[���#	���Iٓ N�u@H���q`�	�&2ӆG�d�����C�{W�5�B�h�SI�xq;mR	��J��+�s�y��g�O��q�iώTL��i���`��x�O� ��~춬F���0�u��g} �Hc1{���_���on1�������Y Ȩ8ߙ�
����֏F�F�$� ���\�e�������D��������ޙh�ûNPM����>�C����Z�}Z�iryRp3Ӕ�F�D!R�]v���k���-7`d��3���������/EI9�)�%�#GC16lm��,U�᤺fC�ա�Aֿ~P�9��|�ͻM��&�`@� w�H<��d��z���Dk}���CMs�I��Ya�E��0*=⥰���R����y�z�J��#'R�%aX�l;g�Mk~����5$@dwM�	��I	-b�HZ"w����(�Y��LYf쨡�Ԗ�h�v�ғ膩0e���]D����|���-6 [G@����}��Lλ��cg8t5�+�g�9,����c�24`5��3bN���lz�#���ǁ]c"�Rd���pI.�CY9��K�t�>!�&T,�V�!JԹ}},����9��1`Z����A��T����ٰ�bd�f�<��]�
��	ʨ/կ��ԑ�kbZWd���M�Nƴc��1 T�@���ktqK��%��9҄�K~�&��b�!'8�yd3=��a�^�;Sk����*5�å��:?������+���0r����3���4��:&*5�[*�\ȑ�/LR�%�&��x6q����^dW�@���k������Ԡ�ۣR�}����>*A�֜�CĊL�He��7��c:(�p�'}I�TU�7�Q��IVG� 3�d
M��tuҶ�6�(Cӷ~�w	�,aѧ�6�>�X��N�Ĺ�-;��7y �$�f�[�	�\���᏶��b}1:͢3�0���I�n�AN`u:v3e-fï��\��+��j���Z���GT�d�Z颯J���$�i�N�S�"}�������4�Z�˰�?.���[w��p[�Y�8�S���g(2��:�*{��>�3*d�)4 ���E�ƆdS��	�;6-��v]�v���N�q�W1V	;��TVZ�J�P�1K�@�5�a��/��V������X�ӏ�����f�=�� ��C�8C��ݱ�G����8W�r=P���E�S}�-����#�848r�p�u [6 5��B���ힵ�%9A�˯,����Kn��j���&u|	�hƁl8��K�Θ3����P���i!���y%H�h�GK���|9��o���+��~��w��u���'�=`� 6n%O�9Y�vՅ�R���=�\�1���	���{���}�j���ŧ���|t� b��� _yS;0e�h?�kW�U����������j�@��d*��x,�?�����kv� �z�?V0�wZ���y�	�䎶���#�t�&̤d�0��7�R?��2xU����vm����*��%EϿ��C�)>dx<vq<|C��Uk����*�s���'U�v��b�iS��nd��)1-��+ǳ��B��bH���ދ{^B�ō���ᒚ����t�����l)1��0 -6���J|�\��+��Qn���;�M�~�A!�mBo�P�Cd�΋��ҘC�*t8��λ�vˠ�OǯՅ��}7�?d���t3������S�o��A��ݸpNv���M}U'���$&�������,Ix�leVz�;<�	�z�u�=Ơ8����2��̪@����ʒ3]�����!�g�k��س���Ɲ�q��PG����P0����sgJ���ɕ�n�>
���䁁L�J�w�f`DF�x=+㺋��Y��	��[�R�i����=��Y�)��Գ�!9T�I�^�
���hs���U��c����<*Ũ�-`�[<0�.�����j<Q
.�Eﴺ܄����ꥻ"�*z/�h���~�nդ�P���z�4��؃���q�u������\O�Ŕ��+O��9!��:����VZd�M��S��}qznu�V���p�z��ѕ�������-��+ʞ����A~t��c�c��U��Y��Gz�x��.5��v��p!G�-Jܵ�.S�#K@��<���{M��e2��o�J%v
�"��A��N����~D�~L