XlxV64EB    2d84     cd0�(E�x�U����v֯b��r��J��`�[+N�wV=E�}�(/ށ���9ܞ��ܿ@̲g��>�0Խ�饖��DV�l<��h�de����c�.ٞ3��	N7'�/�V�8��d����1��*��[��A�	�`�2��M��ii���%߅:�\߯���z�4�W+��A�l��)�iQ �z� Zۃ�9M�3]��GP��a��b�V�`�]��h�G�Y��2�h�f���[2L�e��V}�-��
���,����<g9lVh�'c�?� �%�� ^�ү�J �9�9ф�<���]Ǭ�&j*I��݆��l�1�(��\�}n��4����aN�!�NW+��_�T��5TX!�
'>7\��n�u�<~���$�ȝ�-�s|���TB��6��d�d�}�DW-�h(��!�@?)����j�
/�q�:���N2�nE�BH���)�8Ul%����d�,p��C��D����k�	^��ʻD��xe_��
��6֑�pU�.T�~�$������ϴ�Z3h�RɄ=�z?
�\��>�_�L��$S�4��Ob�CP��܅�\m^��k�P��� vޖy^a�TB�.��G	����I�������	]��rH�$�el"j*|���Gd�R��x��r����ny�Ò1-�Ђ���.x�����*�'٥ft|0�qF<v�Y�6�>PxI�5`���%>C�덫�|�*�6N��`��DOjp�I����/.�,H��ثb̽8K\��J,�>���#����Rdi����� Ͻ{>rjr	dAl�\�^]���-�o؍����L����`#��w�``%��@�w�*��&r�4��0<B�q��GGe�6o��ԏ�!E�n�vT5�곕��"�葥�X]�	1�K<���f"Wh�kE$���~�@h�!�@�^'��g���R��n����?0�f� u"�����r��p�U#�&U�k s1j��6��G��m$�h��H�L�A�'� �f�4��?r���%n������I{cQ�]�݊qS>�Nh=�$��������KN�����3�6}t�􉬺���Vx��rO�S,+��-�	=��S\�T⦴L���&���g�sr�CQʓ#Dl)�jM��v�b,�Nh�݅�+"�v2ݨ�4���b�ȅ4;��*�sW��-��:�ĵ���;�mS�#6%�s�Zz����,#�a���d�j��W�������ft�5���M�6+��)��dd��Z�G ��{:���&��u�ֆ:�_�-�zmL��@h�V�f����hh����-*�ԝ˯�:<7#� ��Z�дq��yŗ1�k>��-���r�>H��U���U���&}1�>UD?��J��L"�X�$ц"9�|�n��Lw�č��0Z�7�bԺH����0�|__����H�;�*s����Vm���*l��b��;d �榸�	�Fۀ�(	9���M�h��V�*�* ��vX�$�0.iu�m�|��D���u?�aPEHZ/Q��*����l���=@�>4R�?<@��c"p�rK��/��麦J����R��8ə����M{��+� {f�r�U��x۠�Ik��o���L<>�gYiG�ގ/݅�����_�-�S?�k�
o�^����P�r{Y�Gv���ՒF�.;ܑ��U��z��FY�- �g�
~Z��Ȼ#��̉���z(Z���s����#pY�#�K� ��Djü	�X"�nk�q]�����@����a�_��"�`����cgG�Jڻ��W�^V.āɐ�={��2OH�#���ͼ��l��`��~�Wr+ӆ�;*�t�`�~�Ȃ�lq_��j�c��u�3cGU��/� �G������5|/YP�[��a!1[��`�yg9o#�_�V#LJh�V{�Q����b�aщ0e[� ����Fw_�&8��	 C׊��o9�*��ᣤ���z��$��� �U#�&����	�tG�@�����9�X��T.��>�ru|�7V��u^"��_�w��U"��^P��0x1}��hIH;ș$������������YP>��;�gK�P}Hzx��?*��K	0q�2�Z�/��l��C�ps=��2����E��p��^�&^[k�L�%8�j���Ԁ�4m\H������)�o�EI�a�Z)&`
{���`�	|(��i�I�
"� [8c�q�z�ȕ��xC�Z�u��?���Z� �Rb����;��A�K�pf�~���>�y�G�.n����k�:���;N���z���,G�=RQ3��w��BC��čYzƒAw�ǘH`ĵ�p����+m���'��b�/�}������[�U��)�x/TQ~/�j�� ����B^Vv�W��,��s>�+�!B<ٔ%��s�,���~��̣�+��!���K�e��,���I�fZ��A��"}��|=���6L�U´�]���'��x��J�"���I�������������;	�j]hl�c��.�Ff�řfҕ��)�g~Wo�[�M��<���o���Ֆ�J0Q��� ���t��pM}��x�c(Y���\�ya��r7*-�rǽ2p2�$~�)�䬚]��O��8��x�L��Sv�!�m�'�¨����"��G���d|p���g�F���v;�E1A0��� 'b��G��ڲ��	1�Q2��� �����Y���M�h[RH�G�E9��k������!Xt`� A]w:`R���d7�R��G`غp��`�y"��[���0�w��~�S5�����g�^��2�l��j-M�熖
����L��RP�<Z�!��j��]�n�v8 Ƞ�pW�s�}����k����l5��8D�k�)���v�]�C�pQy1ɧ�u�X�2؇��Ɔ�����՝����4G\��{]A���#���}������}#��Qvf
��Q�M�%$�A��:��d1��.˺w�P�n7T�a���'�_x$b�,��*�i[ߍ��gt�Q�6��s6��C��vҁ�e��0��^����7��@w?������&1`��L����{��6�aE���j��[�Z*f�W�=���	[�3�[��ѭ����bd�o������|�%��E
�Q���S�x�0o�xO�M��u�_�]�w�M�s_s����C��@�)��U���g<�