XlxV64EB    8a39    1c30���+��~	fD�W�8����/{��Z��xX� !��SaEp��T���#���d��|K�њ�4*��8a�r�����������+z��� �+-�#%�v��r��f��R]f�L����|U2�[�	#��(ߘ�h��F�6xG`!-���9%%_�gBln.@6'������Eo�ٚ�u�l���dq��lX��=z#��#��03p���^x�+����m+���X�u俤�Y�c.s�����{��0��W�X�L;½�Ǔ��
��{v^RmsaB+ץ�L�EL��+�C���"�R_��/��`H�_�+��gyce´E���I�	�h�~~�+Z1Ln�q[��G�����΀��S��r�s��qu���s�0�br2�)�u,�-N�Y9-�'�siO�JN@��]>K��A�>YQ.�r�X4z:��=���SG�s����J���Ux�<���+.-�	)n���6m����R  �Л��s�ϔ��j/pLd�0�ȁO }v���$� �E �4�h �ꏻ<}{Z4ocϏ-Er��t g���6�� �p�c4VY1�^�O �#���E��w��߹D�WZ�bO��e����MN����.Kvp4(��jFE�,��U�2Q��:��L5�?���+�-<�LDT��cea���3��RA�|�\��\j&����r��ѼfȢ�tX��]O��/: ��X����xL�=%�9�L[J����D�F���-�HJF�t�פ:���m��!x����
���g�೘Yrm۰5�k�!T���!%���mu�3fg���;^���9Ģ0u7�R��q��%��/ P��	vE6��uX6�o�I��D�n�3~�v��^r~R/p���x�^�y��
}00�7ԏ�ks�1���/�d�'�/ͬe薥�و�{WD��Kq]�ۼ\؏�-bN&�
=�j�D$��(.��׌����EŘ��4���nƵވI�#?���c��'�9] �MKE&"�M\|u�r�\��g��8�'�aP��Ѝp%Ӻ�@��Vߐ)0[u+z��3��ɀ!�n����M�|��H�$�
JB
���l{c���Ο���3�.ǔ�:�S�x�n�����-g�V�3�Fy���ѳ�e��)�؃g��S�ب.���$K�Zڦ�;b�����s�<��8���r���&�(��T��T_�D��jE�ʑӔ晵<0�� X�����wet����sz|��QC�*U�����_^�m�uP5\}<E"Ao�Q���B�d���/+ܸB_D{@�CNk�SjC=�X��9>�A�oOZ�9I��a��q��|��' z5ҷ�W����F�}�EKf��ģ�~�xy,�?��x����u��R��Hss�=$�]+ ���E��87C�`�JuVe/�+�{��X}�8�쨝�6��daDCN��fD���_t!�Ο~U~��dE���׹�"N�HT�X@�蹖�[�IQ��=_�π=���x��M`����}0���r���]L�2��$@���ЩK��9cM2���z'��*̖A� x4u�e�XYS����n{���'��V"؋,����{\p�M�(�7��GIs���`�e���>�5E�y�,��{*��H0���*�hHAw+��&ڴ�4��+��r�-g�)�� j�3�z�'���[̯g"l�%����k��.o��TB�݅j�yU���՚�8>	r	��b��/�3|�󫱗��xP"�q�i�ł�>����fd�@���k��l(� ;�\ީ�'�Kx��M
pZtV(\˿�E���U.��(����ȑ�
���Y�C�gy�B'�9� ���u����mP��,�݊.�A��<5I���^�a+�R���Hܷ�x����m�#�TG��;�؂\�|�Ґ>O��(y��^i	�g-$�]�,oA���n����=֛��]
ܓ�!��sW��u��G\n�e,���1��7��mE�
@N�GdCDW��|���/��	_S}�X�B��Ї<S6=��x�X�-	Xߝ�l��^D���7;�����i+�����\|���_ߡ|�y0��=������ȟ#��,#�eX�����ǋ`}0����튝.�,�KZ��ob���B�!��3�X{.",�O�<͙����\shM�/��|����~�>t짭iV�'xs�����K�#�� Z�����/��{
�4
�����S.����!���ʨ`��T����uҢa�T3���|�����bH2P���1���M���(4M��$<I�r	Z@
��H��33`׍���)#�[�:{1�.�Ĺ*Q@�6�l��d��Թq����#��L%�Huf!�����;���Riu�U �O"ķ�u,��aV���|Ҍ�1m,R$ؑ=Q�^�����1Sc<�9�۰�?6�ĺ7,�t�S��k��M�EC�p^QbPc�B�)]���r���nErI����G�����"�1ud�ݾ���|�Oj[;Z���b�����G���v��(���U��~�
с�s����.�<���)���>�����i�#tp��D0�N����6���-'
q�&7GM�ѳ|n���w/GՁ�����l[L���e���/X�[���c��t.x��$^��+uy����m#��t:Buҏ��6��G'8��g���&�]} Z�0J-���"޲�N�H6�Zùj_M�&�w0����`��ꭦU㺋���.�8���x���ކ��^h5I��f1��?s�a �c�.�����n�MS'|g��.b\��ř���Ǽ�'���~�Gu��(��K�����g�ވ>�2�sk�:Rͽ�[���A7+���J��6�|�]�W��7��p��B��Ev<$���\�r:]{�Y�e��@��9J&�1�������Q�����ϺaS��5_c��HwwְAvQ�E����	�r?S�daj�4�x.͔���1���?}�,6S�Ň������o��!�nި(����Ţ̢�k 0>J�i�2��	��4�r���*�WM֠�����ܥ+�Lq���_J����ɡ��!����k}��Ī�J=�.&��kn c|S}�禶j�^�䤂�x�">^S 9 x�Uy#VL@Nߢ�H�C��� ��M����\�ѥ����?Ȋ��L�ɀ2��hf6e��^
�/g�.t�
�Kٙ[[�+@�v��������� *����x�[��8*v�� �z��8�-*� ���Ɔ�tpe���C4�Q����@�2�E8<*�f�Ý�����j���!��#��k,͏]��<-0WP|2�I�.V�_BN$
�	� �!���(�y��)`e��mrWn`��m��;-��;td G�Q<
��L���Yr"���N�6�ˋ=> �~㞫��e  ��@@�8�|�n+�"���1����"(f�-��������)�Sg�\�W�aw�$E��]8�h���RR�7ۑ5����iFű�c �Y��)V0�>�߅���2�ߋ���59�
лZ���,��aw�Yny��1L� _@����j���&)�2����̳;n`7�\��i����[����j������Qn�Z�5/�qVf��F'T�Y���眎YbW�6�Y�@���ʢ@k������^5{7[�_ّ���яr2�믚7Hb=���U�kE���v�9{�0x&���[)�֕[�d��b�wԸ��uk��%��p�R��ʩ�s٢��Ķez��eFꓐ+��]�՜F]4��Е���/�Ь��ݜ�$%Xi���0<��q������q �X<`�F�:���f�w�� �4N�v��W����b�i`�'��R�ψ���k��zU�e�N�R�v_�� Ή�_^�.�X��ͅ@�S-.�gǣ���p+�CXR�rߋ��*r��f������995B��LR_��F~q�}Kp� ��^�)P�`p5���x�c�aq����mA���L�n�>0�x(r��%��2�HÖ�06B{�"kh��[�-Jq��1��@�
/y�]ʭ0u�%��������m��X�i��8�+��Sf4@�*�d!�{Ό,�(�7Di���Fn-w��t�������D�yL��Q(��|];0�S�Vt�ډ��Ț\��/�bp$��M�e:��u3f�c](1{9���x1��Ĕ7�[6|,��f�ޫr'93���T��iT��{*|BO����L�m]�S��F���7A�� �$�m��`�)Y�+����nKيd(�?�sEx�ǘDԫ�uB�̚
˷~Oz�r�%D��	:�f`�Q���}�>""?/z/�+F����In��fN��	נ^�i�5n���^&5;�S�,�Â'�g��x��ϑ�l�L�ܠw1�V/�d��Y~:�kR�ќ�0�� �Ɣ�ՊBk��S�r���y�A�a�'�<��H��]h�ReZ�M�)��fx���9�bs��
H��Sө>���
� �ض#�ﭶ���m�+�����?�f/��j��Ǐ�X�p Z�Ym*��y �q�~������$��l�8���
_U�m��tj��+��4��1�w~�f�Q��A#&z�N�ej�<�x^>r�E�eB�P�>A��Q��c����BE�0�'c�Z��|��:��͉a�����u&����P��ȼOJ ��{O���_�j�Sʼ�/�C���z�H��|{�� E����[��
-�68�2~���ت����J X��)G��w��?�Fn@��Ŵ��9�c	��ՋC����� gB���,�Z0�N���*}�]pf�.x�?�b,��/3��3�Xz8T�{$@�l��S���T�-���6���:����jr�$!�)Z�⽤��`æmB�ׯI���vJ\Q���'�:�l�(ҒA�>��>(��
Z�
z�㷧*�DE�z`h2�/��;w<�#6��9u��:��H������w�y-����Q�k�����bG!c`�k4�R��(*���OGa���o0.]?�%F�hL�d��\����|���:�{c�.�������\L�Dp0��TM�����k 
�-e�Y��%�*F�O�C��n[�}���^L	�����v{s��c�0�V�����c��L�L@l����T�nsKޭ���!�L���c�{b<��Ԍ���e��p�:��j��� ^L�>�a�t��|��m�?�SJ�a5��e�tgو�t�Q���c����\Bs��)$/Ca�J\cs<U�EL����������{����n�mLҜl��]�'	�_޴f�������aUF%�Q�D�WӮh6�q��}Z�eD,`Z�C��!)w�.z@9c�>�S��[��,�]��ƿ_2�6A��%�����Km8����^�W�_��>B��*�Q�����I8��[ܘ����[a�o!D�mק,ޡV����L~�H��L}�F��1��h2��I�'��Rq�Y}k+�&e��[�����Mk*���y껲A��mfD�o�z�� ���t� ��kP��)�l}��u�e��D�?e'����o~z܂ Jq"�yx)�3B/i���vB8�1�=r�"�k�)�N t�����X�*,N�M�	�r ���L����nn��nVC��gl�V9ԁYh7޶kբ�k?�/���ۈ�y��Rg�=v�!��ڜ�����𑆜'��jWWA�����h�]Q(�C[6 �M��2��v�ϖ%(���f��?�+S�bp��H�?��a��	ZF${C�ń����������atfW���l�4�G/����Q�-�f�|]�]�H� �B���i,n�#Zu>�gڃsv�(UW?U��ʩ��fS*�K��mK *L�-%���FR�����cru��V+ j�J�;�%o�AΡk�l��L�>F
�6���O9e�������%�F�BP�ũb�w�I��>	&��4_���J�td5��.�������[�Y�=�$?�9c� ��&�7��z�.SSc��ز��<��{3��ct7J3�n=d+�"��/�G��{��t-ʍP�[1�w�e���	lϛ_Q|=�}!OA�¾���'��pW?
��Q'K�����Kd��ccT���7Kc��6�Yڮ�GV(������RM�n�G$6�#��f-���옑�ewF
΍����Â���3o׻�g���@r�'��h+R�X�����Q�����u�q�!��&d��[2�I��Ae���v�@�)K]`���م��h�X���:q�B�'��S&7t�r���uDe�@B�@S�s�*��\�H�k7������=`�_�ir�WqL}��q5���Ts������0�6����E��D�s#��;#�i��w�R}��Rc�������E�4��ce�������;���*1Y��%2��g��f����g���nH�u�F�'ij�z2UJ�������۬v��<�Ş^Z����c���Z/���@�Fp3��& m=a(e��wds��y�Pޯ����`��q̕�HӨ-�������%E���e�i؃J���
I�4��X�{v��q5�s��$RZ9�(��}��%d��h�.��x�D�e���h�f$� V-j��9�]�,�+� �j�iD����#=BM�S���|h�b�t���*��ـSΨ��S�$o����������
����������x�E<�U{�|��9"�HC�%��u��#���H7C$���2�)�Q#ӕ�;uB�o�t�����xZ�U��5�mq��J��$��X�h���r�1������Uk�#�͋_1�}>��mY�|������I	�!2��g���9���`��sz�A��'#c}݇.с#W�@ 
[L�b�7�Uۍ�!6LD��տ�RKt�V�u��<`_�����,1O�W"�nW�^� R(�ks�!�b$�o�sD}V��&�M%�^{mғ��s㟲Iu��공�k6$*���\�� ;��HP*�ĕ�R�^�kX×�f?�zoz
���gƯX���tQu����⳻�	;C�H�hv�A<�Ơu��ɫ�߂	]�5;�A�e�#���ayO���