XlxV64EB    fa00    2220�!g&g}�蘃K�3��lS|	���c?��:m����\�bUt@�ǈ�L*¶�ٞM�L���1���#&,��S2��Ï�0:�)�=�݇%X���=�?>�T�ӆg�eʑq�1uB�ï'��M���k���S�$6ō�i�l~��,�gl���;Jh p;J8�Ւ|��!X_��
	������>9���q�˝b_ �|�]�j%x",��I�pL�6��$M�-���v�KU5���t�,�zJ�:¶|»��Z�5/@��=����3��S�+��?�e$�y�ݕ^����9��ȮK*4*�n}��5`������1��,/�P�� %QutF&<H���*C	"���ް��1�c5�rh���l�^t2ӁŻ�[p!/�Í�'��y��}"�t�6�3K�!���Y�@�92{���L!N쪣@C��q��Viu~������}87Qc,6��VP�3�E���v�D8+�5������P�15cb�]�a�	���G�����P���6�͚�֗����$%j=`7��V�.J,�vI3/|7-�l�Z��ۼ��rc��Vt%�7���J���Wt��8{4ɲ�i�A�R��/j(��ˈdh��0h�����ZU4zc��aX��&n�I?��,�����ͷ�2���c��i^&��Z��c(�a����C�V&�6}1��T����$|�mC^�#ΔP��wHNf���2����[����9�/m��
\�V)G��;��"h��b�4�z�xK�C���\��*V)K�"1�)ت�Ng�D"�I������0��)�%���[�Bs�g:���8�X��u��?��v؟��m	M%�i�	�ry�Q���;��
��*��$�.Ԅ
k�ր!(��o�ݱ�`��[.��߃8�NOs���|Z���Y��F�~���%�v[L=��ڿ;�)���	&]�4�W�QxPdn??����!�A�Y���u}Nύ,��Ō!3=v��(���l�Ԍ�	��B|��n����
b.��j� )�g��^(J���¥���SoC�l�&f	�8���W5�4hĻ 6`����Pe��t)0%�Sa�v��A�r�����
]�]<�������!◧#��^�������0��T�������u�!*��Y�4�r�@У���ؽ-�H�Z�іS�uw���z��I�L�Mn;'�u�?|P}�/�e>���>�$�D"Ҥ�ui�������ˁ��e\�� b�:U���,O���g����^�,z���O2��{�O-Kh�|�oM�L�J	#�b䖹�o:��Gi9��eۇ�GS]}ӛ��H㟫�t���({�2A�ܧɌ��
wpB��l=�4��\�����RB��a�N�� ~�Vgmf�r�an��Ίr�{X��e���j�mSa����h�>[�$"e�����A�o���ͬPVս�<�n��R�5�_28�p-�sŖn��د��z�R�o����Ȓ��ܐ[N�~
f���)U �/�ҷ/�Y~m���~�G�&�eUf�I�򛶱J+p
�,ld�E?:wu��u:E%X��3,b9]�m���q�kw�ȑ�4d��������Qz>���#���7�7h���6�G�S<�Z�׷O]/�FQ�:Qq,sy��������,W[~�.Գ����u�r�)p�:J�z=�����cB�r��h�����v�{6� *X��O���Z��!D)�L����V�pA�[2�	�ʗ���G<R�S�g�ll�vV���YGߧQ���ﻗ ��a,*��4��1y˿|� D�"Y�cL�يC�rz�)�p�_�w�� (j��(T-�������F���U�ޔ�N���������ubj���:uxp�
%,Ì:�@�G/4/bE��n�>y$�o'�I�?+�T��=)�}��������AV�H�.5�W�\'�9j��!2H�v�ED�������6L�᪈a��VIT� $��0��T�c}u��W��A�b��x�+��2�h�=gԪA�����Y��+a�~�O��Y8.a4�ߍ�܈�,���b�i�t�H虔����"(�����C�����`|� �,�v�E�`�}u���툜�1��ߊ$x��"Y���qiS��.�S���0w{�� �zD�\�פEqn��u09G
���n(�M	�֟�M���H��xEWB�Be�ܯ��pWcoЦO����p Q�(�S�v�PfG�r�$FBЁJD���0��U`J��M�K���G�yS��biK"����!�w�Iʅ���ӵ�Kɦ<�}ZӌH�,R��53�%��"�u��OD����*���q�t0�ed�km�ӊ{̇�-6�}Q��Uv�P�N[N��U16�} �eȔԟ��s옹����������Q��oy��>.�Es4R�o�$�n��:��0�`�:�$�gl��=L��u���ǥ��]�Ȃ%RG4h&�B#���O�k�ö@&�F�°�(�,��N"��m1U�9J�Y���$��E�W��(b�k�#wT�R��>2��M���Y�?�o��S$��ii������F̯h��������WNxS��E��Z-�㛓�*��c�7�m�UZn��0T��g��_��:bh�|�<6.ښ�	�>��}�<o
���!oV����T�*}��E�_1��=ҵV?����Y�m#�U ��Gߙx����X,��@8a�^И/��9$��2��1���ѐ������ހ(#i��L�Τ�E4�fzK����:^Ъ�I6GKG��Lj���Y{ꙺ�,�jЖ�l	 �����=�4���v��o�x�N)h�ٗ�I}��c,	�XJ����
���j3ZT���C
��&~��tJ:.my�6Q��M� �TO ��l�"�J�t�O:P5B��r��#춗\�UwIJ1�O:�;SLq:���T��a�Jޠ�A��ؐ���ePrT���0���:����)����D�x\���0��ZY)h���*a4!ϧUR���W�H�u ���==}���H�Ѵ��"7����zb�_�(�H�X�����WP'��&��8�G���n�&��[Cm-'r�؛b��cZ��������T��7��_F+T���.�q��s�Z�覅�]Jf�q��|�8\�H�<4�&?#u�>�yz`�v�jRn�فU�C׌���O1�_d�j�`��&��:4S��X���"/Z���t�ܜ���l��>��J��^��e�#*��ޕ�l��
�B,�t���:T��s��g�.�]F��S�􆂿������v [���&Sa��¹�8!��3x�~����X=T�࢔�ݠ�_T��:��ӣ=��eo���]��՘-e���	M�ۋ姽"qބJ�����GjF{��6��ګ�GL�N�XU:�4b��g�t�Os" �wx���V���&�Id%K��ĉ)��qc����~ö�=��+
��Ł�J������)td���a>�ޮ��DC�b��e[Fས��E=ô�!���>���?�qL|yO�b�����̐|D~�Ef*�{;�꿂7�4��4fk��_�U���d�R�n�kڈ}=���uzS�
u,�X�1�EFV�Q�9A#z�&l[��t�4FI�.G2��"8W�mDt{��S��Պ��s�
p ��5�:���7�e�vYS���C�ދ8�_ƵN$��</[H�o�~p`�0�=_����G ������$S�BT>l�\*��y�<[�_�}����%��J,��,�I
o�ƀ������Vx&{���Gٿ�cθЁ^�$VM��Ch����i�$��H����F!�DC$�v{����UYD��MK��������|_ҹ�B�����Z�7�q���&J
��I׏ּV�a&�v�)�zP�,�-�1E0�a�L�9A�fx`� Dͅ�9:Ɯt���?��u���ɉ�2`'c�U�m�Hf?]�L�Y�\f?��s�6�nޫ@���O�^
=�˪��O��/���%k6ϿX�DtR֙#3��7����>�[�y�m���y�˰�տ����t[���G�a�צ-����
aQY���o�	�~�De�߹@!~�6����Z3�TS��eE������	>Q�/�K,��{r���_d5��^��}�]�2^�� UC��:�m6f �ȀA�h� �SN�=j�xf��OX|>� �H�#A텫��I6m ֛W�gG�+.-���G�#�����
����I��/�X�:q�_%�	��8��8��ֈ�d����ߠSn[����3�5�QY|�S���vx���gz�(�/�)c��2\~A�ǥݒ�����2z���b��0v����t�|�Wb"N�yY���	X�죓����mz�[3�؅kq�7�A����Ȏ�qDzcp�KHP���f)��I�)����\�/�+t����yn'�eXϥ%�`V�F�9PИY�,	��	f�lE�z!�wJ(�M�����낉�=�Qq���L+�:��i�x����;��R�C'���[���m[h�._|~�)6-�M��׆>Pn�H�O��
�����FX�j�{�
zF~����2Z�.Q�`y�
,pD���ص�A������
@}&���������8x�$�T���"�p>w@����l���T`m��1���)�ʄ-�}��פ���W,-�.�����bpdF� �T� �Vοve~��c˔��!7h���V�Zh�m��Y�c���Ur��=$<#!:��l�LB�53�8Bsn�̿��.r]���^�y��ihw:��I�.�y�<��s�\�0�DoE�]�N���`�e��)0�XaG���_�8Բ[BDڹS���T��2�l�-��t��v�6�5L\�=Ή�I��ڋk�}~b�^�uG��v=&�@�(����.Ѐ��.�կ\gO�$8e�u
�� Y�Z� F����R��>����AK6@�8Y)��*�_�L��pc�����4���u�gW ��@5�� -�y�=��ޒ9A�z�_*L��]�8B[t�Zk��FC�6pbn%�:e��+��*�T�W�1�4f�)wb�+��s����I��j)AYGs��y���<̨E���ȵ����r�x�P���5&˃�S���ǙӰhL��Q��]�K�� �L�y��k��Q#�fd�m1J��`�!�e#�ji��`��l^�o�[�n���L�]����K\@�v�i��F>�p�7j�s�{ud�����K���;��/\��b��b����s+i?�]�ɚ\��b�sS��@�P(�����(���s��$3�o��E��X�m�J҈�8������lH�);�n�ڦ�r�^ő�Z��顰��/��y�k�ST��7�KX�J�uU�_��$�M�ߓ�Ac���+W���I��l�(O����"?1�ǲ�Ot7u�H"��m��'���Zy>�0wr�OO�J�2%�$6�N�\
z��K{78��6�vZ_� ����k��<;~���	W�sj�ĝP�i�
�,d��YDI��u�?H;���x���Ms��e��`a�Ov&�J��<R�����zna�J��m��\�t]L�s��Z�ҕ�����*r�XZ���$;��W}jB�={:h�.�m�A��~N�5�2�����޽�a��8e�Ś�_�e�f���	�᭗$��E��jL�z�l˃K8��\L?�����_�"�̡H���Vmig�u=��>������Ĉ9n�L���%�E~?<Y���p�k֦�T�ٙt1]w��`DrM���*O�#�c{H�5��뎒z���L�bs�I�H^�v�|{H'j�Y3z��G�i7�?��b��Ϗ���"y&K�7_*ܙu!3TW����]����R&k��cʮ�����z{Z1�Χ�<a����͑�u �;D�]�����	ΫviR��7������S)��(���0ֻ�6�1��w]�m�9�!hH��^?IqEH�C���᳍��s�*���̾N/�"��'�	�+LW�on�GvqL�#����D�n��6v�\˚h+>�<�U�T=~C��VeT�s���ⱦ�o���f����3)���M��2�jԕ�=��sxNlnB^��4N��"#H�gtO~n��ót��9g@J�PnX��w�0KF����yҊ��U7zT��kV�1����6�(����-���~�]{  OW��7�$�O��uj'z?��јθ�(��ȋ��Yh4��M��<��W�v��q˅Ծ�WE�Z,.sP�W�F\�}����<�ˮ��eث#򆞴{v#�e������#�t�͟ඁ��9b��-�C���ᐛ�o�#�@�G��3+���"Ż��	L�9�UEkcX�6Ol�s�6h/�(��>����2�؎X �W0
Ey9!:'&?>�(��p��'�׺Ɍ\z�t�^dh�@~@��60c�q���
�� V�d1X.���Y&�l������99K�<N�>b�-�=-Cb��|�k7C��Mi��w筠#�	N�~��w&���}�A!��3�R�#ؼ#�#��s������0�atQV�Ht09_1�_Nԝ���G�E���5���H+@4����BZ
�'4������-n����)5b"�ޱb	m+:{��?��Ukg�&��S���=�1MV_n�/�B���"�d�ͤ��4+�S]�5pX���s�������a�G#�O��k6�"H$��xT�c8Y���̡~������-	�>��qV���LW��cy����
����1��Y���R�@����6��y2%��o2���+Ug,'���;��(/��B��F��xu�E��='(o���#Y���9�zx�D,������*7UWY�)���`-�XW��=��"bd�ŝ�_�q�|�v_��?��L���s(a��'~�{��d]("T��M�dխ(E�K5�l�;-+ёDҠ�U��0�v�#���@��J�20r��n��@1w���$�М�B���V����!�U��D����Y�H@G�&����������*q�8� :0���%7�֝M���޹��/�q��z��50�"������?�Q��ʄ�Vt���+�lv�U����v�uT�#+�%g�~~c A�|L��8q�|	;����z��h��E�uIE���]�gZ?a��"M�{�HnL��pH�7��i�]�@iFQ�~�}�7���?�-a�D�.īC��%$ ��%�n�e0 ��\g��[��S	a�����<�`��[Ċ�o��P��\>6V��;xn��5cC1�;+�qW����bB��&G��d���Ǖs����Nx��H׍����Y�f}-�P+���dA,���<\q9�'"�$����O�%��t�����m��>ڻ'���*Lhm�z�.������4/_T$�&�H6�����Qh#2�,�XU�i�-�1+��YnՋ�z;~�w��	֕���Ҋ5K�����ZU2��A	"6MGL�b�+��h�4�$j�i~i�Q#�� Ɋ���gM�R$�G_�:rs����R�k���>����,���B�~�r�I���1K�2��Z�RS�ٟݡZU��^7e�O������P"t�qV�����S���l��5�to��h��wA��%���|��vGK�)��>�`�+.1]E��S|j�n����ـ��h?��M*��t��0���Y����H�w�7,��v�;��LxN�7����)݅��2K��sF��P�=f6nS��Ԕ������������Y.�C��y9CXJ�Ɩ"2��K�;	��#nf�q����X;.�������Z���Y��%�X� ��܂(&�Q�O�X]�1��<���=f�lS=k(0�����Υ��Vp�8D�I��T�O���f%e���g�{I1]S¢��x=�_b�^�-ΞX������r�OA���F�Nk?���Ҍԡ����E��ǔ�l�~ؽ�B�L�QU_qH�6���끦-��x}��EP�V:xӄ�iP��3���3�P�r΋��5T�@��;3�ͲbdC���̼hK'.���X,q�a��s��Z���'�Y�r��I��5|t�~hy�홻��L�ݮ�-76��=�W��>I��q�F���Ț\X+|�b5��/������m�e(�w�Ur�1B����i��ˈɀŕ�^�J��f����=QEW��!�Oj��<��z6�?����ɤ:��R�����G�k�Z銺�o�	�tj�EOtTsʣq�9��9b%k_+�_����)�p�ww� b��
9L�:&1I]�{ݛ����u8<�*�E���O��q�b�0���b�8+�w	
������J]�/b���f��B-k��F9Ix_~����=�m�*X��UXRg���
h����^�$}�j#�UJ*�}��0���4'"Y���\K�"Tu��t�EC�]��^UH%Tӄ�	�C�5\��x����Z6��x���^lRO�G��cd�y��Z�G���(��=�1I�j������!Ѧ�s�*K�"�;���e��(�5t_`_�y� �Y�4|�-��pH ��#ۚ���|XlxV64EB    6cd7     770�8�GP�^+��X�4�(P��*�2�	Z���ч��.��weV�і@���:)n�h9z��=C�0HSAT���(zW�U��~��buHk5�|��e�WE����=�B0���c�2�dפ֩�Qq�����)A�.�s�u�d��_Uu������۾���Y�>j�Pac��+�����n��^�S$$���9���5f��=F''�Trzˍd�0�E�!XK>�j����\5��y�ε��idV��,>�� ���i��*{<��B�kx��;���y�o'��,;f�'$��E�M_�����b֙�h�(�$�f�r,S�Gh8?i�G��6���k��#����6�U"�����7a�?L�9(���2U*>M�����5�ƨJ�a$��72
V>�Kq���'���Df��J�Y�Z��qlDӚt^m^��gY�-�yH�CJ�P����;&�'@#��jB�����q�"����<dc�>�l��%s GB��ؼ�Ȫe����N���˫��w�o�*']��*4�8��7���P�+�=^�\����D%�� 3�v\�����B!�?���h����l�^��(w�������֒)�E�#n���M=˝���[=�{�rNA{���D�
ʻ�tڔɇ���n���O�z��D�< {���6{tC��0�X�W���QET��(�&d�fn� �$�b�JS����:mI0a��8��`7P�}n�r�ӯw@���;t�+M7K$!M�%��-�:�U5���P���*�+6�$>ًҸ�.(�L(�{M^���N�R�j�*���ޯ�s�Ku<�A0IϕՀ� Y"J�j�-�Umj�x�殽�1�5`�N�!����FH���:�U{9d"[x�τ�{�2J�\���t��u����	�k�@�M<x�>��ݴ��={�A�_���V���.�����S'
��OQ�Mw��Mrj���S������ �!�TK����G�L���`��t���ˑ6W��q��u�{������ă~
�[��:�o(��}O�6�0q5}^��	9O|#Q>���{3*�$�B�W��Q*��,I�Y��:�:z�le3�>g�v���n�j��FxsB�J��E`��0��`-�Q��"A��F�}T�P޸q�ئ�k���PN[�!G��X"���
��`��	g���s���g$�ī��C���A���E(=t��9��i!��
|����ևҊ�"s�R*T�QU�"ʿrK<��#U��	9��� �b���B��u`�\�Ż@�\�V%���
A;7�aq�%Ҍ�obs�qQ&{rE,҃hwq��.�i熇�[�0�P;�AB��=�78��e���3�$t@���<Go�/��4D�
�M�0�֚��̚0��Bg ��I���:֩�8���7i�'��F�����YRj���xƒ�<�t[k�,���md3��m9��d-kf\��Ǣi)��p?u;����R�}��"��VF%���?+���� "P%��P�Dw�����[hS����*��a�������e=�*�.��h,��s-{�A�T����[#:6!ط�f���$�[ds��cAEn-&>U
�J��tMx����p�u{&N3�����ݫ��I�\CČ �ɩ/z��=E�^�9ͧ�,���M��-�����>���'�D�`����+(�A\�:L[-�Y�X'/if*�U~�I�H���x#��$Ɔ�S�����(���G�ON>�֧��U3a��0�Q��q�����������vx�"�������:8� �� qoH�T�|87�j�M������Y�-g-�eᏲ��H2�\�|� g�qK��p�-����]