XlxV64EB    6eec    19f0H>�J��QƜ��f�rlb��܍��pG�@�y�Ӄ�+�%X�1z奺~�
�� ezV�nKQ���6�����HR@�(@/A�;�w�.$r����sێ�~-)��*�ߤ H[x/��ܦr2��Z�R��O����r�I�.5����)?��'6��R����?�7�����������yY~�5�3Γ[��b��x��(�����e�9d�50IB��K�I:���$��~T�J;��}�J|�N�s�I��N=��O���
;�`k��׋���|^�!�;�(�-�J�а
F�&Ĉ���Ɲ�P�-�l��K�g����⡷9~�ɼ��;�^�O������~��U$y������FG��r8�
 )�_!�٢Vx4�IGj���7�>����,�:0�QV'���9�7�֜M��!o���t���,�0ࣄ�Qh�}`��L�]1駾����<gn�7O>F���K?Vl��((_���@���>p�|�x)K'gzy39W69@���]�H�٬�:>lT�w��bB��u^�F��s��t�<��Ig��#?lޜ�Y��I�!Z/sP�Z��=�ˠ��Ԇ/�B8��򶂟��qQ���%R���z���U~}=��~q}�
z�TD12�&�lV/����"0�=r��<��H7��<I{G�A蝪b����`���fi���o`����e\8� W�Q�6ش6�yycwT�<b�(��c��b�}�Wȱ�����/uA�#�4�����+xՑ���I�30��s[�S����No������Ʀ�1�맩��)��s�O0�W���E{wPg葹\��id1iu&��=)C� -�V��7n�{p4��uŋ/����� �+q4�)t��6i�ԞB�v��i(�E�o;|���/ܰrr3��.N��6�U�o0���x�4It��tT~����2sl5?���9EzAM�L(����4	(ɭ�X8n�"w���UWIyH̔1�!��]�Ru\]^`�D���뷼�+�]�;PW�.:3p/�raa��mĬ�����SM�������V��_�*݀�'��N�����1�Ꝡ��O� N)D� �4-�GG��;�b� t�����6���c��v���/;��km�yL�xEs��ό��RT'���� k<�����Gyӵ$?2!��:M�b�W�"��%s�����.��Z��ɤ���Q�$!jErOHhu�/�lL�<=z2>j������n+��|/m<Q@�R�B�*jP��B95�.���O.��xq�f�9f�=[XΌ&���� �����P���{B�B�Y��QiK�3X���e�����	��N�i��Pm��� I��#�E'v?�}�<�w��ɦ��="S�
���6����;�+�/�{?h�#��P|��̌%��4� ��l�a�8��[�E1�E�騔�	���*T#��� ���X�o����Z���gT�\0�4R ���n�?ܚv���C�0��i��^g�|@")�&���PҲa�j�YY��	�O]4�S��h`���wU�y�M<D�<����7��!��!Z�����%?�тz'�Z=��?�#Iw�O�ԘhVЇs&yV��[o�[/�Gz��*E�Z�@�EuS�Y����2'��(t������Ȼ0���Ҧ���J?��H��Ju}_��ໞKE���.��;��/Z��e~C���{�aK�����i��/x
��^��d�LM"��e�x��{�O�>�m	�T���}�+䚋B���Gx)��>k���5]n�R��`�I=��3�����'Ӿ�E��@SC��\�֬����J[֡�p/b`0gۿ~3Q�v����������' <�iEg%=P9� Z�W��W��ySvЅ�e= g��Z�Wh�� ��Y>@�y�_Wۢ�V���|�c��F-�`(}|K�Æ�=�J���c0�ge��|)?�;��uU�AJ{���LV~�<q1�o�����wՓ�a	o�YL���5�W��D��z��<�_ª�>��j��������ҁX�ּ�Ϯ|n�?�pB��q�ߘ��4 ��F"�~����A�@���p*Zk��,�)���LGR[�R%�~�U�֮p�&E*;
6�W¹�38{2K�cD��CO.��"������d.�r��*�P��]7� 5HGN�uѮ���t��k����3���S�_WA;��V��+;�s��~6������<�]܏���p�p4�"�j��d��FL�gdbO5�m&��՗u$mΡ�]k,��)u��mW�$�#��&v"m�E(yl��S:V���H��AN/Ɖ	�8.��������R=�\��N�8�kc���ty����̑%]���q�%��i�E��[#t�MCe���KK��L��;�x:&;�����KZ�!�{���ȩ&(MzZ��*��Cē�O�����a"�!%��=����)���BC@)�J��~��F&3xx_������rm�i�|�ٕ�r;$O��Km{�Ģ{;�T�U!�!^��&�:j_ ����"�]!��d�ۣŀ�$�e�;�s���{pS�(��n�W-��9���D�{og>�h�� nUa �vu��-��H<{ܹ�,�Pǭx:��}G3��w�V"�z�v�a`�?&}��#H~�z&�1F^B�-��옮����X��T��C� ��EM�}�y���2�j�]�Ü���R^Js�'��Rh^�1�]D�����J:r��5��c���Y��z��u�s�Vȕ���YDK��民��9��=A��m�5_�e��g����H�o��0����jY����V�d}��ek��=�	��̬~&���(	�ZOeM�����X��Q}Y�l;6�l��O��E�`,b5wi��������"w=�c`�����V���*JAJ]���e�߷j}�Y
�rRo���E3rN����~�@�D�
�qI�ر�	z�ior�+�͊e�;T������9_.�Y����m�3�H/�e�Xk��>���0(7��Ƨ�+a���Ъ�D����g��Z�`ȍ�|p�r*� t�"fT�`?���L܃�=#@�\�k�%�R_3��E4�U������[����^��˕��2!H�̵��9�`�nb=�籠Ux�%��.�+#"b��F�<��RP&��Wߪ�t���>\�n�V�\��!��ߩ����Ґ4�� �b�n?�5~7==�H�.Q�����oL���%�;Y�Å���5������jx}�c�T~Ĥ� ��m~Q���ݮ�0�D-����T��?v7��\�V��7��u�,�����jR������K(g�i��ޯJW�>�� �O��"֖�U:�	�9����"Lx.1z�'�+yP6~��������|9��umV�N�PRFg]��Tď��!�)��tL��} ������~�۳��cu>��)Z�D�4�.%tR����M9���^�>�Lvɰ9�E���JFL�Aw;hU�`3�"��cÝ#l!�uD�O�Μ7z���k��{���.�@:%��}���@ꌴ�������\l#�����g��;��$U���`�B&O�6�p@{��K�EpU��V�EY?"�-hU��R�旓�x����v.�,�Մ����/��1��[<�$����NK�{��Y��L�}���^�<|�����7�'���l���j&�B��ID ���E!!�"���yb�kj�1�>S�1��i0m�Fw ��Ւ�;��J��V�f��"�%�,�٤���\�a�$�����ƼdIQ����8I�u6���rg��_��C��h>?�P������E����
s5768i]�x�⑽&���p�V�x8��;�Q͔ڒ����'*�����iQ��jg�����ϼ�Cb�r���8���������^�|j�i�RW�Y� ^�_o�&���zGd��x���
,��\s�FQ���2�#���6ҽ��C����kH���=���e鹷�����5����~43&�=[����F:�U���[�!��%S��l3Y�X������{��fa�r�!�Dŵ=�2�)9P5�@	��������Rl%�:���A�W ?��ʸZSR�f|,���S�������$���O���P���;��P�;�020[!�6gy��3y2��0�a�*vA���޳�o�-`��ϵ�>/����ʖM,΄,P�����MZ�iTB(J�F=,%F~Yd
ץf��)Z�ǊI�O���?$�����Ԭ� ,��cQ�Q����_u��3�.|c＀�KK�κ�XpA��X��݆�v N����X��	a鶾ৼGSp�c��b�&|d��l H��T!K���9BZ����xQǦ���4��K�@�b��1�a�e��	�5L��F>��GjTv���`��n���]�њ�P*/�]����J>@̵=M\)[��y��9����������b�� �6��ܠ��l��&S�
�W?Z
uy�<�"�����c��[��p�'�|gq��$V��
t|����U��*��W�Q������j���-�V�Z�� [I�]c���p�\%0�$��wǻ���IY���{�e+�OFS���q�@���5��p�j�P���,s���!��gt<�0a.@�%�?�WT�8��'����������l���
�/�>n�#�_��V]��h(�J5�dK�QTQ�;�Q�-����1�֜�IҊ�ftFu"�������0�"5��m8_���&���s�z�CY��~��l" �q�m@�0IK��N�GQ�g��ӷ��Q�z�:X\��5K�3�^U�4M��{H���KB�-��7̉�k�k�w�l.��)����bL��'Z5�hu���D�����/d��J�~�?b}SG�k��~�� ��6?��;�Cta.�c��L��{ ��8��nB܉Ժ�.H3R	���5�J. #A�����w�Ka�L��S y<�E�H�5Blh���Z=��?p��k�Q�����e>��r�	1�~����0���Ji���N�@��_;�����uc��A�k�9�j2��m�(܃M�N~���ڱ\�� /VB��ڶ$j�V~y"2���b��Q�O��X�\e�!���+��^zw;8�~pxO����ƥ:RX���ü�CΦ�|�FS7��23�CM��uP\r	{b��"C��w{�f�㱎\.�+���8��'��f��� �]�E����΀��-w9є�,�/�N� Mj���3�R��?�e3��~)��XA�4��Ɛ����ߙ+��iE��ld^Uo��U�"�U2�?Iw��'СY�2��v�	��X���\#Q|1+�e 6ָ/�<�e'����lkV��:��Fj��A[&����D��P8��0�a������،g/�\>��:]"�᫛s�yT�u$�o�z�BĀh:	���"3�F�d����p��ҫL9������iF����dJ�/�X��ꖈ�	�&f$�·7��;>����M㯪�	OoKk��|� F���HG��N�@my�G�D�Y��Ms�J�BAPy-iOJ����ʈP~̥���I�!p�C��eÑ����y���NK�Zdp4�כC�F;1f����]��$a#�f��~�3��{:[6��} �G�Q���ӗ�oU3b�ؕ�zߛ�����#O��7_g�wG���\5���L�5ʒ���HMr��sO��Ҿ�_��5%6�]]rGO_���uT^�z}b�h	����;�S�E �<%w�ā�S$���@	��Y+5�kƣEaބi�D�����`��=��c��+WĎ �i��	jm�x?+�Ge*�Ѩg2!F���n�q}-ݧtd?K�U|"���	�K/�n�����9p�p��w	�G������9>D2�J�S�mx������\>���З���]�v.��(鲜�Z4��0˿y�jK}�Nn��r�41����>ֱT��{�?	����M1Z���*<	ZkQ��0ʚ�\jd"Eݻ"�&.:��B�.R������!Vr`�������R��=Mq�}�� 0��ǥ���������X��z"@ܓ���&-�|^g�h�++E���ua�s
����J6*a>�VI�w���b�����#��e�����c�n�`��B��߲c-	
xQX����~����k�%Y# >L����3�H���ؙS&8'#\��l�%�ZC�Z\Z���Z��{�7^���:5�⟈n���bQ2�d8r,��W�Z�0M��.`w7����='�jw��4����mz~~��	�����?p!�g޴�,@]���ye�x���n�,����f3�,p>Y*�E��hW��`�I �Q��:4�P�������p�L�b�tXv���߯�8=J�2饴[��$�4}G�	�͈ǩm�l���� L�_B*�,E-�pP��ۻ��S�íF�_�#A��l  ��