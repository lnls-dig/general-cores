XlxV64EB    602b    15c0��sy�mO�f��n�Hm�>��SN8����5�4��Q�[��zI͌�x�1dMn\�0��������R���p�:�(S��F���*R@l���|"a�R뺸T�����I`gX
��|NMwe������p&OJ�r	*��M�R��,�k-��l�b���y��5�A�U9#E�u��v:v�vp�B��e*���a4'��5l_����t�����I w7�4������Vt��)�����  ��Ţ��{wo�RŸ��'�6L63�}�� v�����X���#�F�O��;�{滂� Y����{S��,F��_�H����Y��9�:�m�3~�̈���^ j5PG��l��n{�׫d�������7h�����(k��}��G����	!)�i*�΄�:�۔�x]m���{^޳��	��`N 4;r�:�r���U��S��dDmɓۊ=xiK���N-Cc��R [Kʓ���"���n:ܞ�{�0tf\f�g��aS���7�D�~Fa\����%�B� c�'ޗ\�؈��1���j+t�Q�|��n-nB����ӽ6g?��z��-J���[�����J��=�y��Z��%�`8������j����1DDYSm2>5���DK��B9��'���̫����_&�!L�ʵ�)rZӋ��3��'���+�fi��Hm�U�>$��xks kz�����Zһs���YS$/*A��d[U�<- M��|3����s�P��n�Rr�ɾ�ؿ #q�Vq_q��	*C5ԍ�O~.)�*0�
*?�gi6��v����=�D0of:�~#'pY���
J��4��f0#y�b���M��)_j������=u�=�
ȆA�گ>����NK4���m	�Bq�f���ivY��dho� ��3�]j/��i$���[�v�=���JVnU:7_����uԣ�r�g�@/[���.ob���<cɎ ���VW$=>si4V��f�8<��Fv�/���ӱ���c����G��iW���̣�_M/xd��f^;½�d�6�8�."�0c�\��4r����?R�1N�R���D�W$��"U�����\��h$����珷|��S���Q�)�=�ކq��j���7�s�i;���	c[�X�+�<l�q]xS��Hw+0ܞ@|E�����Y���'{�ʉ߆ʄ�e�ӾIHc%��ݯK������Hԙ�sV��{-V ��YZ���J�]"�K��	�1+ғu!&���������RL[A�������\"Q6�Ϥ{�0?�Q�H�h�c	��X��j�x\7�ú� �*�̻��-]i�G=L�R��!��ßæ�#2����	����Mj�1��ru��"!`W�}4�
�h��)!ZZ�(ʷE����d���Q0�8���	P�>+�#���ڬ�Č5WHN�A7H	�|�����=��*n���YdR8���I��PB�L�(Վz�H�H�C���`���QoCG����H�S�K���̼��-����)�Dn����%A���wu_s�~�&�V�<��L�A#2�Ɏ�P[�כ�e�'޽-�p�\�K��]V��G;���J���@�w#��)�b/���Wwc�����o�d�2�J@ �[�K�s7�X���SM�
�[�iI� ���i�o"P;EݕI�t�!���Mu�̓��F�m�ο���(��� �R�s&r�� �I5ݣ�����x}?L��J����b��▃m�n�3��ÝH�y���(�%��7��� �C�������wn��ߍ᭿�3֍��$�Wb='ׂ��'	1���t��-�QEخ�ƺ�]Gx�J?=[�$UNNa#������0�*�\E��dL�E�k,C��S��Ce�/S�d;��;OZ*�L~WY�VP՝)Oƒ��n�u�QN7�B�]���4\����f ${�ċs�g*r[����v����^�ӕDX�i���G�����ԄJ"W�B��f�2E���m�5 $`�s���2�ʇ�U���9���?-���mEJ8�0��V�5��d[��G�|�5�!cn�
�[L��=EJM
cF@�3oo��I)�_�Dj�S�
H���B���%��e�q��
~ &�K�9����1���|<i^>��[*�y����߉���*�kӥx7u䄇绉��pn5�o���U��h��6MS�E'$����%'$�Jd�^^ȪE6��2p)�� tK��el[r��>�i
�5��4��aV��Zf�KO$/��U�pxל�T�m��0҆'���k1���I�� ۳��t8�4���GWk<��c��@:"Pf���k��u��I�%oq/85��q[�i�b�7p�6����z�	������g�vZ�ڝ\X;^'�Cs��Ȉ�4ܬ�V�}Nt�gx<<�_���� I\��V�sx(�oY_𗪄$ރ51���X���G򊩔S%ZEGSaY�9y\Pmy$�@�ɛtV��<��:�Y�5-�Ka�P��N��O�)��2���oY�/��J:��H�C.UL1��|��G��� �q���?��NEl[a���� D�b-�ve ��}�|����G���/��̱��%����د��f W�L[v+�k���u�'�S�҂�Q(�&e�	��݈.�BOmvG�_��$��]�j�</vT���k����{-�5p���y��5�<yQ��"˕LT����ʱr-X��J���59f�~[`���b����8q�j}AM�i�%�)�'`�+��Y����
�����vI����ս�g�,�\�6�A��&v��W�o��+�x���k.n�I��"�J��ǫ/���jӘ-�_ǈ��U&�|�����8w�c	���;���cvk�w}(���L�b��S%]�9?��sɫ�:���魯�t�_<�R�I��h��Ӗ�tY�}W�珟Y�N�H0���ͫ�o� ���I�X���r�&ԏu�R��g�)9�~�N�灮��٭���c�'��^3G�ۛ+� �=*'�a�fRU&�0���5��d���hL���'�z�&��/�z���c�o`�C;ÃQ��=�8'�s��"���o
����C�1�A�i$����&ڼJ���玱�gO8��%b����۲�u����A/�k}Q��7�6��twa�����W��n��nnS���q��#K��K�Iұ�<�0 �zi����"�uH�z_�i'�nC�U���?��*	j�U�C]����Z��Q^4�
�*%�ѬxK�ϡm]�	9C5Ămi�j��n�V�4���~��N*�� ҫa��O�,�͸�BXv՗�+ ��L�q�l�n��T��Hٕ:�v�6b�7&�"�J�A�:�`�s�-�Q�p����!�H�{��y����s}jU?�A��Z�#nw$F�Jx	̇5ӧ��7RG��jX�&�-��[�G�b���E(���°F��@���m�thSV$><���9QP��*ͭ5No �k�3)bؐ�`�z��I�k�}f�M�8� *�:| ��,�J8�;.nVڑ�8$1H"��������:I�2O1�߉����y�6Mr��_��3��c���p	Oe)E/7PDVa�sn(#���Uպ��>�u/]�y��B�9���q���J�? (5�a���Cj�y�z��i�+��!���@���g�GtcFj~S�����
�g�柖b�L�ޭ�a�CJC5�z��a!�硜���� 1Ѯ�|���b1�W�@�\����dA�̳�g���%J�)�[Qp�Ԣ:4��7^=h��t�xm�ւ��*|�d>9�N����ar�vEy����߮@�T�9�8'|E�'�/���lj��������0Ҥ�A�� ݗIwz~MI����6L1i�]�Mc-HbE��[?V`�4�j��fr�;j� �!��F$'��r+���B�K��!|{ƞ�@�W.�}#�Rٿ-��	?�?�q�(����)Y$x:�R^Ho�!Y,�Cz'�K!���+>��
݂�z���\�zds�´��$�~�گW�>B]���@���Z��+�/C^ab��r� �Q-	]��Pc#5��tp}������%�,l��\q&�O�Q�Z��RqyX�\�`U�4��$�}�l�_�eJ���[���G�P��	3"�bzqA�~��6�2ߜ�ąqF�.*��no���xN�_F���?������H�CnhF���*}��TH���;�ʉs�{���f���E)2�O�$m�a�ˣ�.���D"���=�|vK��g�uVY��hX���"��XW��K�c��Ut�W����{���P@�a��Lc�|���n+�E���C��=�ҁF@	�!N�Q�;�dMh���ӈ@@�vd���3��5��#�R��=q8���NZ����Ro�1��<cWw���$y��މvзk�`Ey�%�o�МH?e
�e�R	�!K}��Ѝ!P���&�'j�]���e�|��̀�]ܥ�C!;l��yï�Qzf�� ���Ǝk9.JLE��[w�7��!>�`�j68 QkՆ4�π3�C�a~�B��J��b���\.;!3!�G��65�oo0Uϙ|��=�c�j#�S��E�����ѓ�ↄߓ��92����J�Pp�`���ҩ���{�#Z4����M%�׉�H
T;���he�&�j�6��X�Um�6��侜��ވa��Y�&v�d�j��ВX��m�"��s3oeQ$� $���G�b%9�t7;���e�!�|�!$H�Ҥ��6��%����������X|X����ϻ1�7U�s�$"���Hף���=��w��C�]�F��J�)0R�E!%�$	D9���|�����{��z,t�F,�����b�Ӝ�tș���n���}JV��EN�>tA�W�y�Bt&�r�h�ܔ��Zda�����+�J3�3�s<W�}�!U*���J����!�1����>s��r
���{~�ƒ��@7�0�z�~B.3����j�wQXǕ�sh.�=�b�������eϟT�\}�m8��*$���C����u�Ԁ؏���1A:�s��!2^��-��|��S1\����b���2nn�.�஦����qB����*��x��5�d+��Z���GTռ^�Ó���z��H��x,��(�-��� �3��L�^4}e�8u��!F %�!e�Wi(b��j �HN3�@疌��cF(R'<�蔐��Q�eS�`L�%�� �5�$U�a*����i��'Sa��"`�Cn�J�%�n�{ewu����<.��-�C�O�IlB�~w����^im�ǝLw����Z{; l��	|�p'm���;����+��$��Gm7����g�$�<:�Ӧ1h����R^�;۠o �0Jj{�\gW��Ay��β_��u#���p����@�c�X��E�(yߗ�r�(���3�*Λ���r퀤#�Yt���2Yݕ�\