XlxV64EB    4684    1090xR{8�c�'����v�:��I�bS`������.��c9���2$5#��r[�t��VG���uKs|���`&-�I�:��@�ģ0$��h�Om;}��=K�� �[y�/X�_��	�)A0�|�7���a�8�&�7�z�Mq�/�r���^�
c���X�����٫c@O��?�@Q�rXL0d����Ί�"(�`��U������~��u�)��P��u5��	��>5N�8/�I�Y�!PU��#b�v�nP�T���� �HI�m[:7YNT:q���!�]�]��۟�@K�N�7���ۙ�о��)qq����I@$���^Ö�y�H�w�F�����!s�G{����=�>��-¯�?�U���d-܆-ҌL�oAN�!�j)�B7ã�\�<?/��uR�8�Y7��7���-؜攓�٥b�5����׷�����J.�j��N��R�b��m(.vp^�	�n?��2u�����݆�da9�*��>о9^.��ч�B���O��=��
1���i�q�ny,�o�����+2G�ٲ�8�6S�˂{��e��#^�#��+�O�zɫ��LkrN[waG�&k��H�گt��K�'y�b��@�"%7N��}�#�\��̮�� �$��ez����q��s$���+��R�V|Ѽ�y�25��Z7R�V���9D�=��c<���'-~�R��o������*29_A�����!���`@���x���O��5!\�y� 3�K�qfz�6QmЮ��Q�tΩ���C��{���v	v�b)c/���(��"	�o~��A�/@�p�]R��Qj�� �`ZT��^��.q_k�Ӆ�.7P4t�sH��+`���O����]���F	�g��W��ngM��-9���G�bm�5���(�׸��[�e�X�;4�P�&s�w���`-�?BbH�*;~�����>���[�F4P�L���6���I����fLR��ޯ��5��O��F��פ��F�~����3ȱ�B��jJ�F�KJ��I��Y[Ĥx�\��I�T,�e?^|4�4c2��z�2D�Dt��>�����2M�ϻ�K��!�Zf~L3<]�j�p_�p=$5`*��'A��YAA<3�������"����d��oiHg/�Yp�瘽�H)�o���z�\I*�r9bz��8��e�U�?��p!G	F�v,���Ev�
�M0$Y5�n�.�3�V�
�rAv);T�
v+!��P��0y��/��5��&r��nTQt9`�>��N/��q^��5J��Þ��n���p��vT;[���ӯFv�@�����i�OBF�M������سc���~�������#p1,DL+ܝ/g�~Op\[�A5D��uI��땘�Q��f�ט���肮��
�8�:!e
�nja��l���~���j�Oܬ_
5�֡8�%L'FW}Q�r�����7f�Hm/�3�����)'V�u�����	��WV�0͏e�|NW.7�<8U�HMp��5Rq�u�}�:p�h'�S�dy����i-+ù�=:@8M"�ݱ�J�)�S�A �ì��¨c"�P���a�x0�EE^�XW_:�%�1Q��T�1��w1���9��Ύ�������|��H�@'Eh.�ل�W6��8�_|bz�U�"F�ð��J���g�]?lX3��l	z�0��V,^�E�j��E@�s��"�^� E�;?��FF�Q�Pb�2V�/�?�c�W���P�?o�2����|>���
`=z6�~�͡ŢkAw)���T}��֍$����b�Nv�6�0�dl�ؼN�ӽSU�I0�oU�-��� �1�r��*�/� ��o�Yǲ������x���L��΋�v�a�1��:n���9���Q��#��K5:;�oO�Y��4&��3�ߝ�t�#h�U*�Ѭh0�H,� pn�H�D�����̒9⚧��4��v%~��}�_��т3��RJ��i�P=��J�m���$��P�^0�1�k@�[
&R����C_\��_�ߘey�)�3�k�@�k:l����%�U)��!��c���X�y3�!X��C�@�K��ŶẒb�񅄊��ۓ�wn��ة��i������Ø���r@r�lK1HQ?�k�אO=����A  ]���
 ��3���zG�6`��I�C΁�\c���X��J�n�ň�[�1gp�����vt8�ߢsnM���Qu��(բӈĔHiL�Hh���6
	ů��eH�ѕA�rp{U�|�!UF�����Rj�E@��VcO���Lғ	��J�;���2�2�м���H���'!A:��+7N���`�Z]�_�yuS���i�O��=u��Z�5���?��T�������9hp�[�p��سX�-�p���=�hT%t��t���qSx��������n��`÷���L噊J2�y/Q DmE�GMnJ���aa}�}�틐[�2��=Wo���,#s��I��h�Y_�>��t����Z�8��(A���0n��yg�	ϔ��[�"�1��:ֽ[�_,���'.v 1�9�2Ҿ��i<R$����r��+�81��;�1Ґp�!R7�[��Zj.��~l&T/��x�ш�91��G6�H���O;��)�5�Hg�Y�l,<2�����t��.&%�#��:���v��},M�$[q_�{�#�{!��1�mb(�?�jV�ƚ3��uG/�5��'�K7��M�	~���5��I�l� 0xe�N�i,w�2bXb���&����
T䟉���"��fV�i���U��v��]�����\�H�������Z{a���;��[��7N�uP��mD�J+рi���-[#�Eu+4ݽ��5mT�|�7�)J�{j�GƖ������V�%�?;H1u&���"#l&T�J��X�TS����d��V!��w���C���N�C�y&��EyJ��~/Ƚ�[{�pk�y*�c�$��B�o�M��)�����[r��o'��ڙ<�o�����[tך)�"��q��B�{�&!l\Ur^� ��E� W�?�3�l�O`�c~���#���$3񬙂`��g�-��t^1�lj��c+L� �	��<!j��
؅aV���J�3��@^�,t���H6�#v[���溒�9:SUA��`��-��nU�����1+V����b̨���?[��]��6�r{��
����¾AY��oj(���K��=숲|�ZL��O�O2ɫ��F({��.~kD�Y�p����؋�_�&J�[������H� ��0��� �a}��t��e�W��G#oѵD�㊶�v���s��ijJ�� ����C�҅cՆ�� ;jg.��YH��c��\�4� �X��qӧ��}�OVy�Q�3�rp)5l�e19���������\S���
Q)QUB�:TPלW�!*����	d-6S-�ܪ�^�^�.������w�C�2��y%7�/��/�?������̯�L�e�V=ΐ��k�0��_A%��ke˧��=d<��;Cڀj)1j�w��'f|EU��~H�5��d"��zwl�P��xg�~����o�póo+2Jr���M�O��Ag?
��8��rl����%ps�1nk�s\'P%��[��� 7C(춏!W�z��!����Qf���Foوh�c�qQ<U��$�aPi.�1��ʶ�k7��X8 A��?��et�&���~��.�r�jz�Tִ�9��&��|LO5n� 	v�Sa�#_!E�Y6���ʐ*Fso�bWGi�`�돜���?��$s$z��lL�}>8t��D�){U����9�4�u*�-@�+���s�m2�����Y��>ۿ�c��;�bǺ�Nr<니.
 �.C$e�F�����D�\A�-AMP@��ɐE	���^��WE�[$��HĊ4F�LV2�*���Q;9+S�Z(���k��J�҆0�_�'���E��k�,�����E����9(n	.�^H7k�/��	�^�/�{�4�pd'nm��D��q��+�Gv\T��P��{/Y��%\����^���rQk�)�,��[�yU�w��R�{Y؛�q�_�-�u�B��h
�>��r�	Ǚ,������=�a�H5�� p�"��h�����-���������}�a7�x�h��V����5��̑�9����M�[0��*���H�Ͽ-�l����