XlxV64EB    fa00    28a0�
:5�2����f2��宼�Զ��\n���p��Fǃ�}L�xaA	�k%�!�'�����64�V��a���PTL�љ������e�a��p��ʅ)��T�`(jHoUQK}�T�Wa!X۩Y-yR�Q�6}S
��� ܍�2v�.T_�2���Su��0�34⧕��l<7�\4Uʰ��Fm!���r"�ٓ5�P�fQ�/?�P��A�Y'��48*���-8�*ؤ��_q����ĳ
u�f�
�#�tW�	�7��2��8_�@��z�|���ZŀdCjBF��$@6��[o�.��%,��@4�����=�11鸐���<-�ء���v�'�9��x�%��TĊ�m� L���=����^g��bY9�&(���zޘ�L�X����Q>�����1����D�=�A��n�����n�	��������m�=��?r���x���ʹ'(1��B"
.���Y�K��\:�jV���Re|·�D�b���T�}:�L�Y�9*Rj�[�I%��}OY��#s]���hw~!�=��j3~�[2L{5IY��d�D�K��	���է���6�C�ʮ$������AU�1��R��o�$!�<+�Ӏo5�2P����y�=��f]�uV�����QH��9�r��_MUU���sz�zQꦼ&�@�bu�#vL	��<�>D���l����+��*��R*&�_8tsm>�<$+6_@ �.���^��Wb|^�ξ��@�ȹwl������:��{0�P�Ǩ��r���qX� �W����'Q,G�z��^6;v[=(�E���?�m��Rj�'�I(h�}*�RnvD�F��~"Q����L��y�p�fo�;�xK]�r"�������}&�s��\�{x�/�5D:n��[ȗ_�CjxZ�����	}���~����H�7]��������]���ge,`e^ƣ1R�쪹�2���P�G�w�E�N��}B��E�w���u�~f�Ԫ�.�!���<�o>D>�ӑ+8iV8�b4_{�צ	�e��_��ք�w�[��q��3�@�������'�!P2n��
u��7z�3���g���˄�}6=��2;��[��2mP�<tM8�i�/����:�@S���ua&���keK�=0cs�����K�.]��E#W^�ȝ�9������{<�xT*�����Т���ojpF�����x�}S���p��$��\��/�S\{}�m�X������va�n��h�=�����I�%���L����<A���+H��+F����,ifj�����.����X�w��F�m7'�Q�X��;��0��2�}������wv��/��_���4Y|w�-8&�0cJ��i�}�Q��� 2��}�DҒ� 6�wI�GNo��%."A/� ҝ������|
q$a
�3�/��I���O|F��>5'�t$]{�mL�?��a����m�T��[	��Vy����4�T5��}��;ծ�ee W�4,{ 	 ��ʵX4pj(pܡ��^��t�3�{U��:�>A{:tx�]�*�4"�#D�/y�����H
��v�L������%�I�,`~q���ހ:�p#$|<7ͫ?��x�c��x��Ls��Z;��K���V����߱���7�wO�E���tP%H��hyפ��, t�b����/����3�D3���
	�и���W�|��Snda�.m�U�����3h��nz}݉�Ϥx��X(I	�H嫡<o����d���.����B�"�F����2c�^������8���7o��=Q�]���M��])2��_�Yw���)���;-42.W#@���o�7�6@5ie���ޠ(�º�?�r_� �GcT��47��b���!6;�d�m�!x��!�D����HH�)���m�+1*I	�/�)@�+s�c�v�W��C���.�TiR�����ɬgd0j�=H�a
)kgrR�*5�:;!��N/^�;�~�v⡣��X�`�E��w�,f��4�-����j`�3�%inwߝ��|�9r�>�Ӝ|ͼ�ܓR��
�j�
:��K^v��E��}�OU�$��h������{����-葵��!����J�Z���EC�j9�T�O���q���3����u� ����5l���E: sX��j_���Kw�K����l�q�S����4�{�3Bd��C�)0�\&��������El����u����ǒf��Et�	�A���D~���f��!K`�F�e�o��j��9�L�j� �[���2@'��M׺�m|�l߳A�a� SD���p.81����VGD*gP����a�����v����}p� Bo(�p�PwY}�j� ���\-9��	;�?��`ޢN�g-�Y����}}zu1��9VŁ=h���s�cb�*}؉Zd�y��!�Ȱe^e�Nj��Nu�lMp��B��g<Ɩ�<n��-1�;�Q|�ֲã�˖t��1�r~���j9gY�����'���`Pdd��z����nc�X]a̓�&��U��?�\U��]?����q&��[4�a0䚭�[����C�����k�	��y�-�|T��s��Ƃ%5Fp�jC�a��ܧ��pTW�x����"ʫQL����A����t1t��%��g����h�^��.L�iZp�f-ۚE[����,Ն"��n�������MO
?>��&��ebl	��E�W`=+��6C���_{n��O!:b�����F�y]�h!��������Q��kS��j�FE$v~��9�{�n
K�����#�P�5�yyn3�6�KQ$�/�o�`?��&`f��$%����?���:�Nc��.d'�&C�����Ftδ*�=�|��=_Enh��%^tG֡�F[_��!�%��j;��_Vm����"�A_�O+�#��m�d0��tM#j#X��&48`�@���������*E��@+�9&ϛ��gc[}�swۏm�1��:��хg�#��V����qD ���abs�[�&"�{����@5�&���!����o��e�ɾ'�����J*�Z�s<�J�����.�~:G�`U��A�K���^�fw?I�
�P��/�xL�G�$�������,żj�� *�@�b�,��O쟧�n��ٰ�(1|�GS��1��&D�3�r�n��Xbo�\7\^��{wa �H�19�f�V����=��^��!�3�t5�W������Ǒ$�{�0�:�"����uؕJZ�T2�bf�#�q�oכ z���9��;�>\��=Q�e�����p����C7
�6 y�h�Ԧ\G.5W���)�Q��z��[�IYF�\��n�_��\�3�(q��n�ě,�m����U<�Wdp9����̼=>VG�Q�B�m.�)��!\�x{J������]܌_.�}�y���q�v�ʹFDa��XI(�v�
e�v�/�����ĭi��'�c���2+C�6a�2	_�e�.З�����o
��.����h� eVw��,���|��)�0�a�އ��3yx��Z*�׽@~�"�T���ʹ�����k�?�����L��Һ�+�����yW�y�E�z��D�~GL�m�ż�n��={%��&��ɴ'/^�Ԯփ�Ƅ����8:��?gh�s�\y�թG����`���Bay�^�T�=�� �&��2�t�~9Plϓf�6�W�9�+���Y�siX� �p��* N��^͈՝���L.�LEISu��#o�I~�5҂ǿ��R���W�q�M��j��4́���ձ�Ƴ���x�����R왌�_1娽3.&��tӍ�h����6�t����c}*aI��w�]�YF�"mSY"�*��MB=��(Q�+�oHv���[�p��@8��}��
���	ߋr��� /]�^��͵�g~�_1ey����b^��	SX��������k_�'�� n`e�{�D�z�^�Cu��/5��QW$�:!���m o/R�+������WKf��qg�F���G4�e eO��ݷ�Q\��3���0g��ϔ��*��;��E/ryh;��4X���
�N,�0�pQ�M
�&_�C�`�_=Ike��%u�aW��u�Y'Ʒ��ёs�D�&����&B��|uiT���͜�^� =�m��O���] ȫ��Ե\[[t�/ۓ@PLbu��v�6*9(����D�I��g�@��y �3#cFMn�}3���և��v�rk��<�a�ղ���y����Ӥ�[Ϸ�[�������t��f�� |���vO��=]R[7���z�������]}q[�v��K����@��.��ā|�.k4:)P/��o.��'�Z���U�T	n�Y��8\;��S2Ӱ���O�EN�Ɛ�7r����2�07��{��m��2丬�5��[�l>z�PB��%n����x~�׉*��gvdR������H�V��䅨�����G��Ԍ!��G!�߽�u`6f_� ]�P@�Rp�Z�fY,�P��빉Z��<5*Ŋ��n�Q��2ָ�+�hu�h�9@cǜ�ڦ��P�;���)i�$ȝ��
o�ҕ���l8�A�K9�Ù�4_�1�/��t(�r#������z���~��-M�x�8�~�.�.���3I��q?NYc�KYI��`��l���\�\�z�I��c}��e�=}����`�h�=�%�I��l��:JJ����k�*����<"�r���wR�)��34W�����!��Xe���R:�ynY>2��F
k���@��ג�����]v86aر� �����qY!��1�b� E�����(Ҙ1c��cѩ���t��sH���Q4Cj�I�~bn0C.��#4�D�#�(˖��l/���a�\f[�>8�}���P��pԘwj�ELg��"A���9����K쭗�%����K�� �|C  i�r�W��O�O@8bǷ">,54�&zն��f��oNhM�\��G'�(׎��2�M�ܺ:.y� ��$�~��M�aq�h>a����Z�~Lez�/��k�o��q���ȇ��O����	���f(���J�ʙ2�q
��(�tj��f�yEl(k-�(�.�εMޞ��"���_��;*F��
8ԗ�rی�z�6�ǒt5�Bwl����W`LҔ�H��?2m ,���nvC ۿ���
J����s�]Ο�'� LQ�e`��褌p}�'\c���0ۊ3V��4��/H��d��L��,:��� ��_<h�I����f��O@=v4���Y���:2�J�l�����)eDli�ɯ80�J�k�н�)���DR*�$��o;�pQ2����ܽ4%��������@l����綕��2�v�lR��Ľ+8?���J���,ՅXz\�dW������|sA�98� ��%#\:#����1���1���)��`YУ��`��()�>�Oӹ�dCh�^zzA&��4�~���}*�5#QJ���X�2:F�s�+R�A��������t��Q1�rᔯ��W�Hl]�9�I#��[<��,��>r wVnBy��~�v���mx�i�°���>S<_t!X���=����q�Uě��]6�%{q�'8[Y͚pǢ�/���K��$O��W���q�g���,f���MB<=�4�Tő�c�8�mE-BZ���C��ij�ٝՒ�Kgo��*��hHD'����X�E�-s a�e�Z%�v�O���i��2����%#�C.[��j[�׽�R�i�t���d��	���c��
��x�[V'� <�+Zzԓ�H�V]��VbJ�ߵ׹v<z��A
�uK>GxĎ)(r��$V���MfTYd��&��r�S����/���g��M7�����U�"���7����G������Yv�`ծL�c��o�m9��M����)���o�/&�E��%��%V4�*q����}�I�t��D�Ͳ�/U�Gua�0��U��W̌d2x
����o���L���_/�3�|�5]x�ΪǽM��w��`�dx���ğ� ��s��z*�";����@sCs��d=
ȃ���%�C��y~��y� �R���=���>������J���2u��rb�������@���t��M�2y��G-�$����W-�����@m���0�����'�6�!)ˡ�$T��@2���s0�2 �-��dI���j��}:
�Qhq
��ZO�"�+/��r�pG�Z�Η�J�-��A�e����{���px[�!������w��"N|]��w<m��?.=�\�>�F��
�h�'�����3O(b*�A���9�
p�r9��Ҹ����9�[�끋Qz'�QH�L��M��{��'�h�'�Ut5���0����ܳ
��sK�R�����(0`.�;���͙�X�|~[��7�Ӎ�K.�������p�n<|�9\�)j�s�H�R@��S���7~�0�RS����)���^'/2�Ve�Jc>��A��HlpXX�xi���|tt�'҅[����f�ЁH���4�W
KT��6�+�7�R�Eg9�[BNMp�O�%%����6����J����O��8 .~"�cuB�d���,=�:���{k���x~�қ �Wg��;cNAxϦK�a�Q"����g>L�"��� d���^,�y�\���S���8S,BnK��D�q����5�\���ŁQ��3e�ѹ�kkgv۪LϠ�Қ-��z�V
2?�f��HO9��N0�o���-���չC�:u�f�uf-k`2�
�{bG��1]�����)#�V	�6m�CE+a%�O�����Ʉ	���'&���"��=^�o8��L#qn���<�6�mɃ%��(q�5D4����?tE��J�8R)#hm�H������kJ�A�~I�转�6wuع�Eʉ+��q�|��+�������C�������+M�ruG�)U���H_���5�
�/�8�硉�+[��JJ�1q�1��T?F���U�C4��VƆ?����,����F���Y����HH�0ɓ�@:$Re��������r��®"�F��ձQ<�x��z�NF�X���C?���M��\��l+�V/WT��C�����aĖ�s(�ў�% G��d��!t:,�E�3�0�c�Ϊ2��&L4���j�{������O.}3�j�k]��B��L�9Y�f�q��a����12
���l���zY��G����R�$���c8�b�|�)/�T6�Y�U�o��k�tF,��F��ů�bPq��{=/�P<!����Q˩5�7Q$���Ar]�l���'b�D*��ަC���'�
L��x-!�l�D�f��_��tW��}�,s?N���3!07���,�6���FA�+��}xu�y�"I�Д��g�3��e~׶��~�G����=�vÌ�"7t�&ʾ�P�o�o!�/��:+1�{5�#�*=+�C�@�v����VԌ/:]�"vࡥ�P��vr.�	��w@�{R"<�Ia?�$��_��#�9����Ƥ��/�&��6��fd��.�7`;�4���j�,ER�me
�Z���-�i��L��)x��R�v��o4T�mG�w��NP�,0ZJ
�m�^�{{����X�7jW����>�sP#/,/�t��!��ΆV�5��=[ �4ԲӾ�p�d,1�a���3J�(�2���W&hHڃd�O�@q:7�L�>���^���!��8�i�+�z�R��0�L�/X\��bi���j�P�#j-���U����L{\�D���(i$5�VNY^�*�8��a��>x�s�jO�,�[�@)v��9T�0������ �2��N-F%� MSI%��zn�;N���o�Ml���=,EM}�c�̹t��'@:���;��"|�-��p*JB�%�Z�Ψ���Շk��ّG����b�ǭWpf��"lo� �,��R&0t��;[%a�
���(uHA���9�s�H�}��5̣i%��U��z�.Ѡ��k��G����T4Î4zeqͩΓ�hr�R�EDr�M���~ͯ8�H�FV�4�o��H��S+s���a����G.#F#����N�
]vu�õ޹���s�����EOM&}����/Z ��o�cN<�QFJ��=إ&�e�7���)/���_a�m�1B�M����Yy��9����c@��O����/;^ٳ�	����ps�&�@��Kz�P�⻭<�G����h��Z<#F\�f����XiU\����%|�oz���1n�	G�gS�p���?���L�QQʎ��wB��Dhq�#6�oB�1��4���&�h�y7z捁=|q|'J�Iж���/Z |��qa��~���+&���
\i���tY�B����G�ARP�~��K���f�?Z=t��l��5�0	iM
�&?�ܯC��TX#�*&�t('M�0�^�qJ��B:Oe\��yy�*��{����G�EOt�N=��j1�$i�G!�ڮ�n?��e�}��ZH!�>.-�t��r+�������B�]j�����u�ؔ��ؐ0*|Y�����}�E��Q�y�P�lq�p�z>�I��G�0�Z��D�W��R{z7D�������.
�\]�DB��8D�O�6�+F��ˆ��i d���ftuK�U�s=��d�C*��
�T����l��?�U��|�Q+�D�[6�|Y*�D�
|sY�z�.���:S��"A����;S�i�����rkya�eC�H�Tw��Θ@(��?ar���cZ~�@�t�Q]���u��ל��@���y3q�0�n�c�us���lB�x` �$C'<�ZQ*qz>jy��}�@�ZLr���s�:5Dڣ;"6���L?sȢLw��ң.ٰ�)U&���ʳy2?��{����:����{ ئi����bj�`sS٫@�]�S��1�&\ٞ�/�Ӣ�y%��}��$�㲐UqE�*b��w���+���L�@	������!����<ٞ��WS�I��cS5)�f�b59IK��F�� �����n\
�kg��о�h#��6	-@gm�"}��b.�� 7�Gn�#y�]�M&��q�7L��u}g�F;c�7g:NQX���~�*y������k�d��^�	$[ꮡ��u�FG�r�� ]����"�=k�GA��f�(�A5Sd�0�\6���6��b4�f�#�����Hܺ��7�R���엨��:䃖��x���cQ�ud�}��ϳ�O4���� ���`q�b����?�y�9���	l��!����ў2}�>�@�el}� ��<���f�L�
��"m#5�d���J3�n�鹢u��c�э�����1�����@�}]�W. ���'��`b����B�Sh��X��z\lBu�_����[5y����&�6}BV?D-?T��/���?1��@�n��X���߾�a��(W'�a��hȗ![�_yA��r�s|�k&����n��u�Mv�'�L$�����ȡ���^�Ԑ:\"&�[��a�Ea3�9���v�?[�C�6?	�^"�������5���!�|��xʥ�
c�,_1/�#$�c��Ӡ�'���b�"��c�4ǰa���u�¹���?����p=?��De*�Յ��_�������k���˃��|�{U��?��1_Uۿ��Jm��
$`�?"M>8�Hv-X�Ċu�E��S�;�%��5p)d����{(�Vz��(P���3�J�=�&bD�j͎}�����e>7�������9^�|�~�{´�dȱ�},�d]�)�.dk����O�$XF1��jv����|�X+�@�I�Lة�J �l����	H^���sD3��3szK�g��YiJ��]<0a�C�oK��K�c��Z�ж��_�	�A*ZO)ŝ�y�"�t��p~ \��%��΁N��&����z���-=�K���=���{:���'�_h�U�?��r���j ۲��>m���"	�ܔ�ȕI��觃B�W��7~$;X쏦�%w֞�<;)>����pW�j�z�|�fz6��i�0�)�W�Z��)���7$Llb��������}n�
�5:^G��YC��2v�_"��vڌw��7�dȳ�,T�N2�Y�qG��P�l�D���"2���R�4�Vwf�r
?І����������x<ȓ$Ͷ��ԏ{pz1����SW*R���/�h>��`
a�[!];�hOUR{�(�Y��c+g�k���Fή���ǆT���.�b(�ŽXlxV64EB     d77     2d0A�4g�z��f����k*��7�l�%�G�����K�C�Q��D%J�uءYZ�$��y7�~W�ʛ��;��{�!��:�7�^]=RS�ڴQn�ء_�?�%@��+���2��t�]`�����v����k_9�^�S!�*�O�c-�L�`١V[v��R�M�Ai�����f?�Y��u�, ]j�A�agL� �������]��%D��v�IH�q��-eNpm���&{/�D L��P�"���,[Q�����
�'$�q]�������FŹǖ�Z�%��{j��;r�hP�:�	��6'�O�Z�\����=��'49Ʈ@4<�xd_j�B]��C@Nm���x�l��QH�\���H�~�6��h�(��:����L�U`i.�!YF��H�Y�Gr�	4CŊ�9�b!%G^�L�IpH7d�@���퀑��G��8��!�tb[��������;��_�:��I]�k@M00Rw~|�X�R\Os�95p*� B�H��F��n�uC\O%��m��W4��x�+�䔲-	�G��@B��$�}��sЇ���j ���C�+�u3���7ڌ'[^w�lXo�(��{����2�,o&��'ҜsF��w(ى_� y��w�w��
!h˷O�XL�6�9*�d?���ԇ��`R��Ft��o-�(K�}�|D��>�C�{��0��g�e���	q��h;V���Q^