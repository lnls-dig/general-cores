XlxV64EB    fa00    28e0���.u��xQ8C���ēt�9m���&dBl@�9�t�;�����J��h#�v�7(�����)"��f^�/VS�<�uf��3������
���p���*�G6�C]H������6�����x�xh��n�����r��J��1��",_$&�gK>�D��?��}C�ߡ��<�tn췯���[tv�N{ "�y.������m�9�gR%É�l��w�h�B����8�j� R}�@�A�n,
�[8ܤI)���Jco���>`�T~"���Ta�M���"B7`^$�!�B9Q�� T�6[{'��O:����܅�GL�Tp@�x�٘�-���E�2VJP�07�˟�9	U����A�6f6uABA;�ޕ1"�`��D��a������x�Xco�
fK��m%X(gW�n��5���'��V'�o��m�Ө�*`0�����pU=O&�=�\��iXB�y�ϽB]xv{@�$�/���f{;?����v�A��y�#��j���}�$���r���N#���\��j���(�� )�1[�!�i3�D3�E�d];�L`YX������xl1DY���yK����?gv��<��l�&�m��Id�c,�����=����n<=nmu�����,]>
�1`��2�Hք�H��[���<�s_��
'cc��u�0D$��!Z�L�g�l�^��5�l� ���O�[��:��V�pEy��g_Jm�����Dl�b��^X#�() �rͱ�ؽZM7���7W}_+�-)�}B�����8xC���wk�����3�Mp��7�l �R�����f����t��C�m��L_�B����(Ύ-��՞�	xUX��B��2�e��ح:;/�_ծ&H�ߣ�5y��/_��*vj���i}��5�-�e@� j�ḛ����LU6=����F2v"o���|6��)�Rv
������C͉��A���5�9j'��=���q�47�GMP�x���t�_ӝmR�kE@�Dū}Ui��TP/+�S`��ca�/����]L�\v��ko��i�(
3G1��o���[ˤ��~9`�E5���S"�*.N,/�IRP{��}�Z+��_�2`�Ss�6��<3W�n�F��XaC8�6_QÏ�{U�v�L�|�iR�
?���zQZ��7������aV�Y �yuc�͊+U�m����c�U��3��7].Yw�i4Yd�e���`���!�f�Q%���d��F���uXM��̒8�>L�@��7�q��N�#N嚟7����O$W�#+�����b�a�$V�Q���s�B7	.�8_ƺ)aI��o�R���`Z��=���V(�{��N�����?����k��?I9`���t& '�Ș�dؿ�z��V��-a���$�]V?((b-���r�Eۃ=0� �F7�O�$%Z|�>��&"�fd^��b�'z�\a�U�\���
��x�3�T��,��Y=��3c�!��	�i��������ow/�/���B�#h���������62��૫�Q+w9]l�N2uE���ý����3�7�BO�[ý]g���]���U������.�2jv�
���$�k����'I��|�)���x	�����DI[�7�d���W��!	F���	'].��2��í�%��|"K5i���g��uP�q%V��:C�9ʺ*�~l��iˀ�SU�C� ��+xY�p�]$39��LO���!��h[L�	178��U��?�������b��!\ɮ��,�������Ilի�C����5c�̬C`���k�[UO���z��` 	�y���rc�fuV�歯d�P�3�6*� E��֮�<�����?]��B�d[}��و�,5V���O_�s�n!���H!���o*�-���G�ǁw	Vӷ���ީXQ�l�����;��s<D��)
����#��!���YU �ĳ���7�K�W-!��9ц���F��m&WV�y˙�_�h��7�*}x��L�F&��J�Q��UX�LO	�\i�0�z�dW�E�ۡ���\6%�^�N&p/9�M�$���B��2%J��Z��pr/┇����O����G3��{>0!-'�Ρ*�	�C�C�Ѫ4���W��� ��ME,T�Qe��b�����Q�A�qNoC��O�π�24َ��Y	lD���'x�-4՞�1"��+�{-y�A{F�v}��$��_����K jt���gQ]���C���]�ML�Z��ȵ+4��p##b��/�0������H��ZR�lA��~eGM���I��y4B=����j���j�m�2�� ��dud�"��h������Z�Z������̔����ǫ�Ԯ�������/(͙p _\�t2���Z%�s�RU��!Ж,���� ��Ǒ����I��{�>�l�u���,ʵRht�3'�^����E]���nը*y� �D�;ܷ�[�t�&I����q{�`�0�U`�MWs��&':��J2PHz&������~ �_� ��w�N�r��n�o�O� �ɚ�;�)�o�4�\�(�t�a o������zR��#�,���(�/5��;�Q�Y��ޫ�:]�����c�����z"���7�#�XRU��\��!Ð� !��}�qXr<�<�� �u��Z�6S���*�2�}����t��Jb��))i��ULr h`,(��z��v��\��.c�5!�Ce���t���ʃ�dN��.�r�g/9��վZ�y����U䬷d�հ���L��N��\�g���S~xq�H��i~�d.I;�	��@�XT	C%��㥤�O��,�h���}�|��l7�gq	$Y	=~���!���:r�����^(�W�/n����>��9���68M��Z� ]t�Ϯ݁���JWG��I
싈��yt<��VZNv��4�H�#�8�H�;�&ݵRx�
��1���ڔ����i�;y<x�L�dDXA�D�P�%`4٬<m�a?����Y5�����X��t���Ҍ��!�X�_jy�b(v�R 4�W?��~ث7e3��;�Q�{�?�:3��[�H���U0�6��n��8S�qL�0ג������$��&n��+.W��sqV���U����	�xY� ��a������v2���e��k*B"���xZ"����M,{�����A�_�sKp�O�̨y
�4��ٰ2H�0j/��a,�D�6���=�.a�-����9� �"R�����;�?��?:�����M�HL�v|��$�`B��u-��P8*'�7��#f{p����f<���h�(��a��k§ˑ������u��{��@%�T�|pv�z�q[*�ٳ�cȉGh�$���y�|O|��)���"1�}l�3�á��AB�w�U�ԛ!�)О�4��;O:cFT���kL�Ex�|�AeC|�4�јĝ%�d�VL�d/�;��Nj���\�g�ćia:��l ������E�$����q���6tq�y�g��38;�F��Ɏ�S�R��G�X�K:�8��
�����ͥK�p'��RֈB+X��m���g\X.W�j\�����ū�ם.�)���.�5���^BE�U���д�`�aT�mz��^G|#����UL&B)v;C��0�:�"�K�S�}�����U�����A�ޝ6هJ��P�W_��(��껳BY�N�����E��:��+��\Ծv��f]PF�q��ߐ��
��~�&æg���@���8�/����"Q�zZKg�(���{��}B�>�x1��w��~Kc����^��J�\,��\6��W��׽��vZ�~f2���JY2�GY1� u�,����h0��Q�@(Vw�x��}�YT[q�yǆ���ɇ2�)�;�o��Ws؉��O�}�Y��A�A�6�·��|hmyG���Y����)}�\lo��LC��H$�T�yG���$y$���fm��g���#��ǯX����Y^h5���$�k(����o1|���b�\
� ���E���ٛ�����|L�bi^�aI"�
����4&��������0�F���,:�ϣZCki_�o�P3w|J
XCC>wҺ�*j�b[m�ye.7τ�>YI��3T�c�xGv�4�~��z��g�B� x#.ן�9p`�s��P|[j�r��(C��G3%��j-���Y2���3��V�m%G��K�U�I�^v�y�m`��Zv$8k�M3�*0$Ys;#��2_!�N�Y8�h�8G20:4vˏ�q:��'�ɚd*�!����޵ �9\[M"��8}/�V�>nIc4�wXW�H�g��)BuJ{���/۽�`6����)aR,�E�j�w��­�Z��'T�4w�wfw,4িm}��tr�1���/�$�
R��2�2q�uD8���zUv��wаMH���]R9ߪ�t�F^���4*�f�P��vB��n��� E>ַ]RG��ش=���M��a�.�g��Gg��쯾),�=Ǟ�WU{�=/��f���?1c�����x���C���d��T�#��Z5>@Vf�VJ�M�8����%�%�x(�R�a%FR�b_A\�l@$Q��34�8�Ay��	q���Nz�7�w����e-�q�0�Hཱ�X����e��n>�Hd�6���y8�&\�M�p}(Rs�d�-�?^ϐP4��(25��%������(����y��	/%��㇗Έ�J��uTx��G��KT��m g���0��d����9d#���?
�u!�� =�>����Ŋ%Suj�?xs��s���J����&4<I�~ݤF�<�K$�Wì
�*J�=������M�A��D��JА��GW�i����B@�z:�Rw�3�"ℭ&-̬��3�T��j��r�hW����]�������[�P�Sг���O�F;�򺽿�����ӈ�j�y����J���W];��\.f:�0]��%x�Tg��~�p�!*5	߉_�����D�+�ļ���j��lcc���,OXf�!X��J�[
;�R {x�����5^���0[������G�	�Ct�ٸ�Rut�y���n�ָ?����ۢ��C.n��8g�/���[eL��A�������'�t�D��BIOf4Z��0'ٙ��ޕj�zr��6�h��M�)�!v��@����-��H�̾�mWt����46ܔ�&sǛ�7Ыǣ�9DĊ�G!�����{��G�s�ѕ�%C1;�/U '����8� �n2)Iw��>��DI�a,ٵvo�5]K9_�-��'��fgXm��؏QW�.�_��C�O1�Q�8��afY�];�.��5H$N�xS�]�p���2�6�:0�C�2���چ�֝/���s��!��Z�O�O�|�l]��v�e?>!����? ��,��Q<��«͌�!jp�ڡ!�B,��׹9��y!�<�A��8���y�D .g1�[��f��>�-�j!�����]�
�|���lN���8�t=`���c�a�Gz@>����Ǳ���W���u���QOmt��^�}��c+JKa�}����m�d���J�5F��XY��[R�vsa���z �j���_�A{;5g�R#-�{D7{].�	�z�jZ/�E0���c���V�`�"�W��)BBu6C��h���=��f��q/�����-����#���{L����.�xM(��۳�b��֞¼_ ��Fm�"-oF|�����Q���]́_��~9����&�K��i� Sb�@w6����U;��7� 4զ/!��k�}�3��i\]&3�+��cp�5Cb��.|�9�ܾ/��) �҂fy$TԸ0-�Y����n�:)+�.�U�/a�"%�U�u��nM�Z�୸�B�K�Ɣ+�o�r~q��F��
�*As�!GU-Uv-���D���8�b�ү�u��NWs�K[g�b�
�)ɿ�6�O����Cn?���>����1�ѭ֎W�Ԫ�sx�' ��وD@�Wo�!a�;2rn�"cٝ�6-
��$]���[i}���������}�����H>�o��E��!���c��@��'K��?x�<K��o��-mBO~���eQO��g���\�f\NlS(��H�7e�Ȃaj�N��>#t�:�'i�y0@/�E�߻8 ����NdvG�I���7GH��J��1?��(�p�w�� �W�P�Mx3��6��Ȼ$�o6@s�wTFW�Ǝ	�0��y�S���+��7g��}��d�G
��*!L�&9w�].�+5�����4��Å�K*�c�������3���@�n$R������#p���s�d��bNe&4Y�;�*�������X�>e׏
�h2J�C�`�ѭ��=�\��<~�%(M�E��Ob��s�ְ$��_ɵN�W�D�Hi|K.���-l�U��ML�͓���ټ��y��E�3h�]`��W�u��'g|=C�p� �*����S;��m����VFł�ʌ�7�#z/"��ï$��H{UvĞV����g��@T���.��*�l/Yн�(�YV��=��U
�9�[���a1�V���a��s;^GT���|��
(���K�{��u44���x)P�J^D�_�(㼆�=K��z(��lRQc�lf��?�i"�]T�qQθ�:��N�x�R��T�'vd8mM�,8y�o���M�A�7θ�	v˻��oF
8�U�(�p��̴���9p���}S�>��:�����s�-���E�ۏ� K�����Ů[� ��J�=:mDKC){����#"lv2�}F 
K�����1_�>�e벍��9�݉��C�%HvH� �,����g����R񪘌��5bd" ��`��vE��o�4ç`�)`|��7�TA|�?�Y*8�_]��y�~N�~�����E^�X��B�	j&WZ��U��2{��'���6G�j��Y�9j��Xs��]�l�4�p�#�e����Q ѯ�F���5�$��#�����Z���jF�W[����ӫ�B��L��*���K�/�?|���O�@��g��X�3ccJ&\tǸ��ėj�=��g���ǒף�*�ѹ��>I9��u0�Sn��/�W��nmg"z���Q���<�FY<�ֆ�����[�=�u$��#\F|�\����2�q�t�#��L�	L
�\v�T��ϑ.z���3�|��n������k���6/q�?��5UnqQܿ^��X2V�#m�r|A=3rsKѥW2\2#{y�Jq�8�������c�D��^��HF�)�.�L��:]��?�����%C�/�� ��
,]�sg.Y��Vrf�˖��EH�L�l7�SH�7Cv��d٫���s�P��*wt��W�a��̈́��6�F��Ws(c-j�����J?��s��4Y�9��Xެd�'h�.ӧ~ħ�T�$�e�C�S���B���y�4���2S����ـG�%n�S�!M�~��k�e�&�r��UCM��-�	kr����X)�X������T;���͚p��$���X���|�����W��\�@��������d�.����հ��y
��.���ڊn?����@��!ou~�q�odA�C��l���E���Z�aw�#�qq0F��5}�)����~���^6��K��[�x>E�i�'#/���[�s�D�s,3��S��"�n�i%��WI��H����.��l�\�F?��_a!7��sn:�B���z��������g��P�!�p�PF#����M�ih�/��}_��Tf�%��F!��o��K6�� v8�%?ɦPB����*}����W���Jk)���g��nR�Jo� A �1����Cap�eifZ6sA��^�	"F��ߣWD�=��|c�
:�h~�6>����Gn���v�\߮.�w�1_�~��PND��ό�tT"�_�Ǣ7W��cQ�͍sʈ��_��/G*�¡��i�sx����O��L)0��/9��jP&��^�?�ڃ�@��B�>4^ڲ��p+����4�^�5!=���ݪh�#S�#�u��rޓ�L���Zۀ��r%1-�K�, 1�c�Ѽ��k>�Ȅ������5l�}g�aEr�e�O���4�X��-�;u�'�%tb���6V��B5�U\ý}n�.��`6'���أ��k�����P�	�ƪ^�v9E|����Oh�����_� �S~��E'��,����h-�~r����5�w��TٝDh�m����?gPT ��E��m��7�9�fIT�R�z�o<"�E*Q�\�h��^����K�ئp�����e��Y-#��v:!��ا�aq�4�R�����X�������I��&'g
��H����\)N7O�E60?X���1q���>h�������DgUW��bt:\L��+�]��:��Y�@���ȀŔ���̕�z��z�pg����53D,x���Hޜ-��H�:�SHd��Ս�o^Lט�	@:���w�����r��g���a��G��S�p|����]��Q���T3��L���Y�}'Șh���H_v�FT\�P�F|�z�1SWSN?�3N~�2�fx��/��G�)5��	��t�$�Y�:~6�#�=���Xߗ���n�
1�v/eՒ.\����VO�)�,�zu�9�$uL}}=�L����+H]�oBg9vϊݒ���<��1�&K)�hJ������*������"��{'m�2��95CZ؋dB����"��5��۩���%�*3=	@�ق���~��_W�3!��o��40�i��E0*�;$�)�@}��]�� �Q`M�[�|�P`|p�i�%���(��Z�9Z޸s�t��_�c���˞z^���8�Bq�_�
��ޙ/F�'��1$zN���Sߑ�f���?��z�~�*�m�I���L�sj4��2���3�[޸�-�1R^�r���r�K�a���D1�T {If�ar��^��7m��Z�i�d����N�Jj#s��K�q�2�(W���n�H����V�-X�,�P3hL+�FF��'�������LD��P�'{蔕mKzeϲ�q��J�& W�\ ��ۯ,X784���:
��b䤕��70"'G��,�1\�~�4E{� ��U��C@hl����,�V��h�ٸ�rQ�d�e<�@A�K�i� k�{°��^�]4�V����m������E.J��W�JXq�_�BZ�Q��"mw;���@_��^;�M���N�$ �Y����/��6��鈒�_m2/طB8�¹�Ëc�o�@L�k�KIa\;|��pLt~{�`��eI���Mt��x����P(�@v���X�rg��sQ�&�Ry���b��8��a�6U 2B_GH+�E�����-jw1R����D	H�kR�yׁ=4-�h���_V(�)�V��%��C�����4�3^�6����b�F��81��J�`�c@ί&�SڵDFֶ�����j��}���G/)y��z��	�	�8�����ʆ3�K;�e��jd!�_�p�v鯽�@5C1�����]� ��**0�U�d�[��M���6L"�(�މi�ٸG�+��_%0`�q�J��ī�kN�9��)�2{)p �-L�%���[�+�(k��X���v�cv)j��>�aU�:�,��Z���1���/(�|U���gh|�k�$fo�j�����"�ɗ���97��%�_���Z����o���Pc0�0�bԾ^���7xR� �L�b�6v(b�&��-ʍ�s��3�Ŗ`���u8�nBKߠ�YT/]�G�-���U8�D�B>a�>�и&KHm���(+Tz�v&M��Ӟ�fA#7��=��`_��E߆�)L
�2?���TXL"@3"L=�{ી���)�7�r�� wf OT��� #�ݨ��Q��%�u�8֓��y|�0��Oh�V�8�]o����LSŒ���K����I�B�/��˔�՝Z����>����bg����F�o8}����՞a�F`���!�"*�e@��.�wGo?�E]|�tS����cE���m[�e�C�o���հuf�`	��@����i�1~��İĄ%�[goVj�1�Izs{j���ք�`P��C[�����!�t� �B7KV���0a���7�D8�Y%bp2�0����l��F�ډ�Uﳲ 4Y��M������D���
�I�gj��$����.�S�U�5*x�ƽ}����M����y+-��E����b��@]E֧�֭�KbMj���R��mn�ig��
n��P��JvÄ�_X@ ��p�Z=�WL���XlxV64EB    fa00    1d80_��m}����Ӵ�@e��d�X����k:3复<9Ck��Υvp�\�yc{��?�k�ez.5���Լ�2:�%��'�|���=�`�׎J,S�sv�3)�w8
>){SĠ��S�)�&P�� �/l�*Quɼ���"&����^䙶ޱ��ф�ݹ8,�Y�ϭ�{Y:���Gi�4VO'A�^7b�ñ��,=��$[��JK�e��}���/1��$_��Ϟ{���� ݯ�v0Km;|�M^O,5���&�����Id�X Q��."B���~�5����4}�e�i���j;p��<�<v���܍� �ɋ���ą�%�h�w���2ީ ��G�w�}��]�����ޟ�1�?�*�b�9�/b�`£�����X3Qs�S���J,�b��}��_-����t�m��qJWJP�ڰ��Ӈ��byT�B�2��O%>��Z����0�8�0/�h:>�	Z�)��?�Bg��D��iKk�X}|����Wqs	g��Wu����zNw�ihʦ]���֚V�N�A-D�C?Q�遬h�p��A��{�ĕ�j8@�k�hɡ��V�M(̋`Is�@ep��|�n"�Av'���m��@Ǣl#��~̅󪪐�7Ζ��X�L������Ė��Yz�C�X���?sU1�@�v=k'��N5�:����L)�����ea�����[KE��Va��4N<U�G���C*^ޫ�ׇ�|�T#'�: �!z�D���3���%e
T���Ȓ���6V+� IM�u��1ht�Mv�O��E��s����ܦ��;��H%y��G�W��Y/��:n�h��!:�ij�(���vs*��u:������¾
J�6)��#�]=�6�pi����SM���V?�Hu8$�Jؒ����o��P����l*�'�Pm��k,޸�@�G�X��)�TL��t$��+s��=ױ{!#��p�Q@�[�E��$�xkK���C����BnTI�42�Oxj:.�Yn�M�r����y�A0� q<��}���<_d�ⱐUF�=��i�4��>DH�S�����	�-3�A�����dM�~�jz�'�-��tΎq����Mx�4�����b��ڋ>���p�C���fu�q�%r��q�f�c^�>��&b}@�{���ȩpnC����!����Ň#���E� 8�keQz ,�h����qr'����$�PLY��i��nc��8=N�c���q�ݿ*�$R���"H	�sn�y�Y/433�!��|�Q�C
�,�,=HIΓ�����w(�k�^�T����ǂn�֮/cH��d!�0�P��Ei#�ф�y��'��������}0�R�Vz�?�G��(�i�
 ~3���������,�B9KzT4v>g�������l�7;΀��s��uN��f*�/���bg����:�
��z�mP�5u�	�Pт��I�������@\ ��[-�Ll�|�m���L�\���fl��P|K��ܒ�O��UY�������Ϛ�\[��`���{H*���!��l\�)��8���r��f-L����>ՊB��v����$�2�X�e6
�����b��A�x?��Ta	߬�e���?'��tF3A7�J�݈2m�#_a*%>2��?0���,-^�	;t���SX�����Vj_�6U��ho�qx����q�H�l�i:�VS�m��!�w1H%�"�.��|>��fss���{~+S�8�_=�7���zD�	8ӄ)�m���+&eСm��|�M�`��������4`�a��N� �䑠�~H�o�>j��CJy�I�1�l&+�Y����L��ctŴ��7=�(�=@,����?����?�i?�xY�5䏸�Ѿ��G|>��*=w��������s���:r/��4��C��Br�RS]ژW�wo:�̯篲���ݠ�]B0�=n{��k�Ց��=e�%}ٱO<Kd�n�B/�WU6�wz�T]�C�)��tV�h�*��)c�,���J����+Fю�o�]�zC���M�2���ia!��I�IզL5W�hZ��'��9�����=��r�@�>��c~"�f��6$3��js6�����q1�9N���� Й)9(IvqVoJu͍I������$
0��A�?�"���E�t?L�`�]Ϳ�����@ ���$ (�M��NVy+M!Iu΀��Aԛ�L��Qj��6�֘�	pw�.'�^�xV��1׻y�M��=�ϵ���0Ӯ��,;��0�*Nџ\�㴺���K74���Մׁ��Q�I�&|
b�4�Ql��I,Zh٢mBqY�hz0�=����a�v��z�@ܤĎ�U"چ�n���'��&'l~��6��N*��pݩ��KO�ՌA�r����Ή �R4��2@��HW�! c�\��Q�w�5�����6���7��۞I3�Pŝ'W㗌���+C�������_��Zk����2TVfs8�r=Q��w
c�r_Cb���W�4�&����C$�ߴ
�]�/�����k"ow��ȯ�z��1yr��˝���X�	R��e�S!G�S����{ik�?�2t��� ?�M}�̧�W&n��{��1_lg�%/Mo���'��[+�����R�J��9��zg3�~.[q�߫�,[�8D�A�O���y���HZ��O=� �/��J���d�r��8�7'��e���M���r�}��S5I=�ș����;k:B ?���;�˾�d�fz�d�k��;)�d�"2"���=q�[2@BT�Q�7�l$F���xf
c{�[�~_#���):�Vf^N��>���Ї��y�(������,�Q�5ɓ�Or$��쬚.�����̎�$L�s�/��Cٌ����F����P{�9�yx�^��Y��3y�g=�Q/�l}����E\	��lI��塁�S Qa�xQkyb��+�����Ӫ�iw�Ҷ�� O���v:>�����T�t�rM^�?5�b6���s#j~����Z��:��0����.I�(
��B��BW���J���<DxʾZ� vs&!\���7=Ӻl���7������U�9��:X�H�ʖ���y�Z�@_��E��}�0�C������\�ƀ!����@���3���՛ğ�WZ�=����CIs��r�h��ΥHÀh�@�"�s��S�gF�n��Z�d�+)gh�0Ǣ�;� ׂ%};R�:�EЈTǃa����ֲBZ{�u㬆���~�'Z�RLO�PT�Nm�y��3g-`6������Zϰ�Oo &����T�L�d��B��"����K �����s��K�(u�li/�r�>��9�z't��QU�v&шG�O�ߡ][�B�j�ɱ��a�I�/*��������X�\���)}�Cr����=�&�g�,�#��L��`
�ϓ/���8U�����MLM.��:*�7HP��Ah�r�qrgL93�a���hJ���ݽ�6��Ob̩�nщQ]ƌNTY4��{O�e�Iu13/�.<� j��4�T�����]iʑ��^���� ����hp2��v�=}�6 0֡���R�C�("<dkK�lP@zБ*�,��-Uj9��N����ZKy���h����F	FT-�6��{�k�	�'c��'�<
�����Q�����!=]�mx?#�.�FY��*q��э$���A$o�%t��1򗖝�8e+��lW��������y5~�b�s!�� 2,���& ��|�]V�3����?��,=�T��<]r�О��4���>{��H�y$�D���*�G���F��EE����U�}w̝�[H���uE��k<�0F����όS�͆�4�2��eZ�)�X�-��7Mn�xT��˴��iMS���������8��GXojyTXzR,��Ox�k[6k�A|�Xۊ�B%�z�V�F'X��1z�H�(R{������sr����/3�����w9��
L��FѪ��A��S:g���n����w���B�e������?�h+��߆`�y�Re�Q�z΀����A1�����^��?��Y�:ُ��zP�]_�)���f��ID�/� ���v	"�%1ZtWBX�:�. 5L-Pwx���o��:+6�o��N��77�.��o=�nc�a�xMG���Q���N�rp����8н 5�0/��>^��"�'b�U�c�)�ͪ�����>B��T�du 3y��?�_T��E�U �#�juI�Z/�v28��;$� *Lx��vA�C�tX�1����\�1-ʇG]����Ґ��S:}5�=� |��+�F��3{�%WCA�yu�2>�_����Q.̣֧�X�����!�YqW1��TT����}q�#Mhj�K�Lf�<��,��H����]̽#����-\�F���Sy���k��`�fǅ�,��!���.?��c#U���(̧4��~;`P-�����Q{��g7!�,NX-P�V$����v6�ITl��/���Dv`!��+zOxt��z�m�� ��C�Z�sp��f���N/�Y�'�����/L��N:q��~�|)��a)�ǲD�r�-L��?PE�*��}q�`���Q��@�7�̠;KFMh�}
��/�3!�8���.�,p!� ���H�7"�R"�QNJ<Nm�e�G��qW���6���k�)2�2�C�t*�ە<�z�,�vQ�$�.&�n��#=޵3Wh�9]W�����X����u�l;�	�� l�Bͬ�{�a�"9d�L�� ��X�M��4��D��p�#1�1�#Ւ�@���i��Phh�9���N`O�KN_rdb*/��&<bV��)Z4��7fD�>+��&i��?���6(,K�rN��|�If��3���y#_s}�M��g���ztBT�b�Z���U�d�?ٰmƣ�g��(q�>�S �Z>��m�!��Y�eo���lo��kQ92hS���a�!�w�^��N��� ��RK8Z��%a�h./o@�7cYAHr� ˙X��*nc.�]��X}<4/iˏ�
[�c}����iTG�5&���ꆒ�?����&!v�NO>�C��I��$5�Ȏ���)<um(���lg�)#���k��l��<�Ӳ <�$� �>Q;�|{qGg$�2�!]G�ҖPS�D�@u��ki(B�x�Np�{�fKFt����F��B�d*ug:ㄓ=q����0Pq������P��cj� �P*"������K1<��_^��ީ���8�0���O�CH���`
�-{%tj���y^ ����946u[�;P�2��l^�K�YYx��0��)8}��γ�i�]ղ�K��u�B���w@Dx����)�ý���4�SL�_�6sN�CiE��\k'�H��Y�dw���U��>�����Ǆ��Ɉ�BYO�e���Iu�hR9.k�������
�l`�i!�d��mr�S����৏$��U�=~�	���$B�;�|lІ�m�zm :���:�o�G�l�惩�-�h�gF5;�I ��fKkH"�V݊��Jǲ��0�ى!��!xَ�-CH�X���,�g��nh�V���Sh�|�_7W&�]�3 űoq��^�抭����4ؔ����"5_� �t�����콦!�Gz��ǈ�q% :j��+��vMəb�4���́�A��u���g(�Gt�,�c�#���%0�
@EH���_k%Yf\�Qu����>D�ʋRb$8�"�t��5�O�<�d�>��1F�� �H6�5�]�8�����ґ32�/V{�'�
8��!2� �+R��n1�Lz��P������tӕ�C/��}Ȳ��+�=�R��G/��������t
��X_��]ϖP��HE$��g��b���)�������4�ʸ�N��=���wc"�;�/x�s���C�j�<+������p8,��L�������(��U��)W��0�&w2~���oX�"��*����wD�Ů/f����M�z�A�六��Eg����<|�UQ�b��cAqI�#�7గ��j?rO/��~��e�U8�E5Z��H��%&���XT�$���E�
1�DP��o;��6�|t�� 좩ѫYVѣ��5ٳ�����ד~����>��5�9[I���jk�����n֙*G�S_m6a>`�8>��xP�1ֆU5 �F��	�jP�1�Bt�W�$a=J'��ҷRz���;�1ORgY�胋Ll�qA���D/#R�Ӭ�[�9<�H��҆�����2��t�l>�f$t������r��������u
�7���n��0��G��#�K�$��<e�^	��4�T }� yt�%�Y��iL�޴[��j&�%a�&j��n
,����V����3�������]�I�����i��_�z@U����h2b���GLR�j: +�\s�y��;.D�Wbn�bȪ��k:(�yYh���(�:T�d�GX�c�� ��Qj��m��9���DȘ٦�w�ۤ�=n�(ͽ�r�9��d.�(/��A���G��#�S�a9��E8pw�G��7�b1A�
�pM
���'���C��~,`ޙ�+���
n�HA�Ġ��f���J��ԫ��&�Y�6[U8)~w�2vq@�q_C;��w'�"*���(~0������dx]�~R3�M̩�S��tyR-t#t� y�H9z)�4�@S~��#=�D��?�8��=4b���k�(t^�tƼK���$gӾ�;��`�'��J3ɪ\�44܋����s��b#Ź����		�2cX�_ONr|I�i7���O��Woa�$Cʎ%���q�6���B`�����,s0���X���!ȑr��<���T?vp�>��	�t�g�,WnΙ���/��
��e�B�w�;���;\�Bu�;��֢R������N+�Ӌ\���$8����k��@����jɸb�̛=�ʄ90�89�x��c�"����1 [:��	 �X"`m�gt0&�� `,a��s��ܑ�zْb+���g�;H�C�����6Eꠏ���}h} �X1%Q�T�d�1��d	��yq�ʵ��T�<|��npdi.}Gڥٮ6^�z+s�U�\ Ԣ	�+ς	���B`b��J��Jwz1nKf����i��5���-<Y{��^s���Dp�0N>��,�r��F�1A�8�1p#		�J�|�CT��.���3b�QZ�j���.AL�,�ç���X.��N��R���M�5�~X}{�D�&ۓ�I[�#��~uY�
� �B��$��6���K��CsD�E2D�Yn&���C���G��_��]33T,Fr��eW��:u8�UNEk̴'�"{mh�5��)o����'J%\�f Vc���!,�7acX?ƹ�=Δ���t�uXlxV64EB    fa00    1e00�u��^j�ø��܊��o������.0G�G̒~֐k�IUJ��<�������W^�ȚR�8���B�*��F���s�_D�r��Z
�I~rjW�{� ���Jr�v�fz��2$��/�H��ׅ(:r	��I�{���-�Lm$}**���S8�N\��2`خ��$���u~�K>�p7���;��!������/�W�x�q�,B�羻!�
B�C�NEW2$s��
�� ��9Â�����
���/sgZ@+���IM��2����e<�Ԉ��!'7����R)�����U'$w.;@�o)莨�6��c�� �f��4���7�>AkqT{�6�Sv1� o���S��:��l1��H@Vgr�,�삠�^b�� l����%h�09V8�J�G&�\��� �s?!�п�A?�si��)�=̘5�(����"E�?G[���m9�,�:I�u�B��J���ݜ�\O7�f�+�9!�4*3U��Ua{ޑE�x��
Q��uԚd!��r��.8x�xԐ��n^��62���|=����L*���*Rz�J5����(�"�K~v>�ȶPpw	�\H6�ȧu�;}:�'(�S����Q��S�~B��g��̿��0f�/���A�j �AC2h"���M��@)>ղ�n�_k�f�9�U2�B_����[���Ob�(w��;U<����B�	��kMrT_wt1����~&���Ӷ�u-[* $����e~�/y�X�x�'X��`pӋy/&@����~}ނg�sm��t�+H�5�󻙎RN M�B�}��X$5s o~��"-�Q��ߎ�^g�&wv=�ѧ ��ix��.�s��w��G�ϳ�銻����4x��O��SK���7

�:�vI�hBP�"�Tj���g���5�%B�R�b�Y�j��ٱ�ɶ�k+�l}� i%vͬ
�uT��k���)��Q�$f��F'�
��F�Q{y�:�:WZz'}�js�WU�Ɇ�?��;ۡZ��N��S+�3��Q`LH�g��4|(�:��Q����=�9���_2VQ��a?��U��ÿ2=�?;S˕�;	FJs�ykR\�$d��|[�ӀVb�V&����[X�����KW*�T�w^U���=��US����3��C��l�_aU���?�@���j��#��F�JTX�4��˼�h_8��������uT�m�u�z��=�:���
K"aX��M��<�sS�㛚��O$_�h��Võ�0D-$7ӹZ��4I1���O�6U������be�͡-b��Kw�B�\�a^;	9�#�����򃹿�4�N���x�4SK.��H|cPN�׵��_~�-5�U���{3�� ȯ��,��~�&
��7�2�N����8ef��R�*s8'1�=7R n�%wt��V�1�(��$x��ϋ���vAG����Xq]�`��{����M�ҁ���B#Ԁ�u,h��n�!�"��ƅ`#��@�h�1GY��6��h���K��"?��D�Wb�Ϝ-�z-^��x��I1}����7D`{ϫ�rԿ�"s�*�w�.�
�=R�'�ZW���X7ը������4��zؓ9�L�oJFR4�*�fo�������l���.�#10��j��D�I�����?� ��i�.Fd����1�S
�b�WK'=���� RnÑ��g��p�:4ʏ��:wh8jBR P#�f.Z ٌ���"4��J3J&�����׻�r�jϤ��2Ȇ}H��Y��u�Ò�@��>)v�T�n�:�KhG'{0�埦�M�Q��l��"�E!�9.��N��~7��_ࡉ�^d�	�V6���,H��4�ɞU͕	0�2K��$޹,j��"l_7�9O �0i�^T+-�<���&w����}V��a��[4É�b��%���3+:� �NH:�5�՜ݨ�s�7x=�>'��+�U��~G��S|���M�[�e?�i��qt�|��h�lL-�[�dx��<l�@��;��r�G�x�v��=w[z._�a��&������lND1�o��Y�Fp�`;�Q+su�\!�1RS�Jj<�ln�K�FВ/�X� ?�EY�k�U:Ժ#�c�w�1�`�!!�ڂa�䩙�ޅ�S+al�/d{�����d�Q����=��<<�dCyܚ�|�����M�mGh�����^��Kn~o�Q�g#|&l^�!�r��(��e���HDR�i-��diCO��;x��t��eN9����@�� ��n(_�"C�M?���45\�Y��S"�K��9�q`���G-��OB$�!��w�>��U;������b�u5�hl`-�#rz)��{�&pb�BX���J>���\Ƽn:7����D_Xo���C4��>cᅺ�/��e�nI5�I��ZH��X+2zJ�So	T}��$A`S�,���;
� DG�Xklk�ηeQ���d�Ƿ�-o7䴂��Z� � l�0晁����s���]L�.ّٚ�<��Q紩 ,M��`�[4-ʜX�ʝ-� �[�����Eυ �w�@�ǣ��0�ج-m�~m��ሎLR¿ �1�7�;�UY�\b���o�nO���+>�c~���EmPw�`�x�xY��,y��VK0�5]��!���P�g�'%�0.�ީf����<����P.��_ [�ngK7Ƚ~�
�TB��\�"p�1X&͂͖v[�14�L��k< +��뉹��b�Y��7�5��l����Mȩ��-s+%8�h"(�n�ݮ���,-�F�JA����F�'(�.��"i\|����@�V�ꇨ~{IJ���|&�;��l�v v�Y ��ƺ6 Z/sV~���{�j������J|�b����$#�;l#)le��= 8�^q��k �$�0�rk����d�3���~�fme�O]/�͂������/�O��<�}d���Ї!$c�x�Yᥞ� P�{��ܷ�)g+(,%0��s�a��`�po٦ߑ��ݗ��w�bhR����TC)������y^ͬ�����@���ķ*s�>4 ��&���%��Y�2�!��U	<
/]���
�|J��£Dm�9V���c-��1�,��FS�+�	D�{t��[l2����A��	�5Wوa2>-V4�����^��z�A��X>"��ɽB��9?.k�����?��!=�Pِ��m'%
 �砮! ��)�g�%��s�:BM�F�N1�c���C�`D��l
�rB˪�ɫ�{�y��'c�~Z�W��	�3*��Ⲑ�����@4���I�BCd&��Vӹ�O���XF)H�������*Z�Y�I��O�!�}�,ݙ����}�Y�W�R	V)����u��V\�ʝ~D�Ѯ�h�S�����%���	�W"���Vq��ֿ�ɥ��t#ہ!��!�lJ(Sjl=�S1�����j����Mw�|����3o���]�'o�t��蟃�����;fV���z��$wW���q�z���O�Ξw�5���1Ls�Ի-]2����p�6_*�[��v'w2�u࠴�'f�����@y��lҭM6ZL�3}V����E$v��a��S�.�[=ʼG���V%�kO�7	u(g���D���P2�jk07�ԬA��}_�&��W35� ��*,�"�E���
��V��?�Ԓ✇��12�$,��꼉�
02
Z�/�dUm�h�'�ͥ�@R^��Mn���̖�
'�-��"Z���Q���xZ��P�c�ѢB��@�{��|PND&��٢��ч� �u5�7��|� ���#{Y�Y�e�r%��#Bt����>RWG9���_3p�_vt��0�V&�%���W�o����]!���5�t'i;}J^m[7�������Q "�6�Ek���PEe+$E}�x)$Xsa'��*9����\6A�p�Pܲ|��wk��"L����&�1�����TY��g�Y2n��-���tM.���A��wo �%'���b�04��ާO	#&g�!��=qD��%��T7o�o&oiؗ�Ũ����D�6˘j}3[�4,��ds{�B�[���e�L��\�TtGk����"���͞���lT}j8�=���W7Pp
m3�@�֭}v���a��14���X���&^�@���b��D,Yn��v�'����8����9*%�,K���y��`,�I�N<�g�Ze>��G
����9�ɭ�lx���(�JM��v�&��]�(~�}�ߊ޶�-H�6'�i��E˫��H�
�xq6��)%��_�SY'�%^U'\�DUF/r�Q���j�}����̣%�f�A��ZG�����<͇�x��P%G�0����Q�Xݭ�p��U��\�yŽ����A��1��&Wo��e��,  [E%�/ӧ��~��]�@̋�L���ࡦ�u߀o�Ř���(�Tܚ������v,o;��}=b�Sg��<���0���UV>� ��]��3�T�%kA�@R���]G���qĜ*�X#Kև��Z�2�H�5d�ֿ�����)pX�s^�L�!`6�*�|Q�=k�@F9�8���[
w����~�@�C�,�����`�hxG�+�5�`�*�Sn>T�U���
#j�[�]g�K�g�\�rfKs�)��ៀ�W�?Kk���f�A5�j�!|��v��K\�L������Oh�V���<�e%e��4ҩ��]+�r�4���7>"�o�J�~r|� �Y#=�����p`���mĝ��UVu\"��;�H�޾���;>������Q�^i��|�]�F"f}*8>��,�'�����;��M�n�XA����!�XL�K�掹4�Z�E,%A�m������eDP�)_p�'���%���B
+�w��g��r0���ڡ�΄���f>�n�q|=}�& ���!�VQO���F�6�EQaB�� ig�~h�Ő޶�L�M�h���ӲD1/W�b��޲8TA��'dv�v�,��=�kp��\.�fL�#2��QO2�I�K|��;07�=r|p����(迉�2k�|��5<�+��W���N��M�ɿYA ��6��*K�."�ʖDok�m�|���Ci���Z���Z%p����jd~j�gw��V'Zc�t�}hUo�1�L�yL�~���<�A�-��٬ׄ/ǅ�Q�6E���ڳ��ܬ���O�@$�˄^�Y�����eQ9G��Y�jd4I��G�ީ��Dm뇝'?����U�p��KX�����@��m5ֈ0�#r.�D�^h�6ǨJ�b����fVm`}²�>m��N��O�Y�8;��G�4jkޱ�IBY���4�py�.SÊ��G����ԿA����!nԃ"�|��F�w���Be�W�G��p���/�2�ôfux��ec��i��وc�S�"��Uҷ�tG�<pNo�u�6ؗ�'LlNR�E��ML��׈I/�)bھ�
�$?5eG0D�-s
�#�ZGt���~ �V ��WBф����t��k>��v�$����=�2\�H��|����1�VI<�^�Y�Tk�MT��HBq����20E�)�  M��d������6<O� �ɰ���H�<'�ȋ��ePP���K�ڿ��cGw�T]oo��,w>��0�x�;d˳�+��V���?���|5H��2�7-�O"su9��w�.�Dug���G�-�\n$����;gm��F�љ�{-U!͢���Ȳe��L ��͕n�U�$8�0ч
|kh�t�=_yEAP�eo���^��g�C��ۦ�wc�3NoD�4�ȱMxm܌�U�-�"7?����B��������W���SQx7�dq�t��_��tq��`�緈��	O�Mv�ԉDH7X��.�l� Lک�U���E~�@���-�����H�]}��c���Y�-��H�x$@�#?h"��r��	�8g�43E�_��Q�Џ}K(,�� H����4��?�K8t��3��sD�2����@�>W�k�)��z�xPf�i�C���+}���6�d�Y�z�D�BS$��I!y&:U�@�kƄ�;T�F���/�LZy��*����V-*-}�ûBlk�[�j��O�f�/�=��G�ά�����M9�'ӊ��$3[���CdQ�I,s���7����WlI H	%�
6ce���c�7����׹�4�S�j�Y}M�S!젽Z��jC���$n7x�K�8ZX҄���al�@Fx5c&m��HM�~h���6��أ�F]�.;�:��c�*����&�����)�~���xPͶ)�T�9HSQ[�
C)�óM��$K��䦿EAj9�|�	��Sǹl~��O�&"6�l��r�Umi
[� ������ǉ��6��/?c��l����kZ���&"[�l�3��`��k�����zjB=y�&���zn��Ͼ�� �??1�Rʫ���B�ҳ�f���Y��R.a�5$aZ��d)��׵J�k>F��te}s ��'h6�ތ��|����`�JώR	�sm��x�0.,3͖�T�8�M9g�|�j{LΌۓ!�\���)�<CXF���L���4���yX4�*�X�Pj\�_	�%=^o	����aZ����[Eb��u�R�ݴ5��)(졛�������K��ժ���Etcw117���p �86<���:�ͤ��cK�WA&�`$c(��k�#w��ac@���0��:0� -$�S�m����i>`5_ǃ�XO�d	0��Y%X����|�Z�
l����$���+��0�%�U6�K9$���uOY@�XLn�
�\ &��ػ�SQ�ȶ���:¼��En�r��d	f���Z�t
g�VdX��`q���ۺ*��7��`-�ٗx_0�z�Ơ��C��-����z�A���哄!���lGx/�!TO[@Km�t$��)�4��4�c
�j+�NO�����%���k�U�j��@�K����[��X�/)�x�(_#=���l��/�gk�1��W�c�y@mA��#@��Q���0� XY=��u��b,61e��� ʗ����h�^�({{Jbc��j~�V�ۋ��u���SPW6�m�]�Q��5����N"��La	��ҽ�R��Ϫ�ć6*�]�du�83�^���7Oت[<���t/����Ǘ|b�e�>��}/���gL���f+�7�ث����1&0̑�-8[.��R6hV�焱X��$]Ȁ""eP
.��E�{ny�6h�MU{|xig�Ll�9�e���$�j��a�oEb��_Uz6�� �= �)\���ۢEcQ)y��ҳ�֛�ݿVp�,�i�6b��;�){�����K}�h[T���2d*��. ,��B���5�]�m�N�BO�f�K����g��6{�=fX�3~l(p]���4t_�����bz��a�w:tw�/&j��֜��f��`߳p�7���NWD2L����. \�� $�F�dQ��	�l�;ZBp�0���DO�?\���;���o?K�fFQ���0.4�J9�ߕg�x�~��&�Pj�mqUx����!���%}
�f4�~/���zÒܰ^��[�����^�?
s�W�{��,}7��
T��'d�]���,�XlxV64EB    b222    14e0�a�#Ѣ�o�,�g�RD�e����~G�\-�I,��.az7nd�-8* ���Q$�Q���D��^C�rJ��� ���<ǥ<�$�C,;�2�:uh���� 	�1��J)
Φ��ݰ�ϖjUy9���i&/��&��(���gsO��S��u�!��22����t�H����W�~����ɍ�ʯO_����	��b����6Gi1G�\	 �Zȝ'M���+��Ձ� 3�Ѐ��'�JZ�f�*��+����0�#�UԡUpS�g\5���k��	�^'!H.�wM�?�a�8�=�އ��4h5�m��#���Dg�X7٭�{8F��C8V-�N]������Z%ޘ�I纡�)y�L��a���<p�:斳:�����d��w��P4���M�r��Nv9��>s%��p�BŦ[.�2��T�`���Bf?Qf�1MiCR�0�4��5k	�\��oosy��}��[�i���z�)���%����y�َ]�b��Q	�ծ������	-�)V�J�B6Z����ۏ����x!fJyUj��rtR�q&de�& �޲��=��(5m���ێ
U�Z�g��W�g���гkY�YU��kS�SJ�h����98����Ǆ��K��{6Oe�-��[�Y�"�����2�OőD���7�Fg'+T�:� ��0=��Z������r��rq.�UL��)F�8J]l���.���89�S��?�5�N�}AۗI�y���
5j���G�]��e�*��l��E��ݫ��k#������3��+�uǻ*.s��B��}$D��gq�����H�Z����?��P@�z@����>�(r�!�؞�CJ���C�����4M����<��夌�s;������5�.��v�_��	�U�^,�`��0����߫42�c�M����~��-9ƣ��������J��Go�T��W,P� L8��qd����1e5��%AdbbQޣ��O�)��c��m]|r{إo)����0,��@�,c�4��#�±Ho�P	++i	<}�P��d ��t�K̳�����MհU���g���Ft������2�����IM������/����h��5�����Wg������2Y�167���E�>SW� �~�i��_�]�!-�{۫�X�K _�	~@��vW����j����b�RQ�7%�2�H����;e��5W�K|LE&�����]!���D1*�q����%i���L��(>L�k�-���
�e{�t��G�+��
*���>>N�L`}>����a#&X?5����5�^��л�1aa^4�)��
������Fw����,��J\`W��H����gN�;xכi	#oI��{�'� A�I����P>��-�t��G5�5ЖKE����.g1�a�]ː-��qI���/ ���0�oߋa"J�`�p#PJㆇ���~O����ʪ�.����������4�����[_C1;��q��¦�5@�, ��TWC��t�9���ƶ��(I޴]]�8�<>y*NƻKוw[�@J��o�^����\�D�`�T��򄴄��$���]lGMt�=��dW搡u�LT�<��z�ϵK����Ѕ�C�:�MY�<0q�Y؁��v�67\^�P�S����1�^�<h��w�Q�fkR�mc�,/�<|9��³[�`}����`/�W�h.�e/9��5K��*dh"��I������3�u��7��������(�O�eCI�p�]A�v��F?�T�H��U�J��%Z�ez���l=���_
�E>���PO������!����X�I=��#'�Ł71P��:pS��.���yo�e],\�0��q�V8������"�Ƥ�-�����S�Uء�,���7�#F=v�UF@���L !`�.��)�?F3�q��"�u/���FeLBPG�F�= ԙ��K;fu�*�h�#l��ͩ�У����D���Ƃt��lt$Vc��v��W���P�lfa���b`�\��L��!p[�~�õ"� ��9P8�m=�QV��.0�$l řn���k<����U�0�z��]	α?���Rw ��4уs��"�d��z������������q	�m-XaLۏ˼�bqQ��mvup5)*O���/�J<�@n�
�1-������@�uz��!��^;�:g��p�R'g��p��u=����g��A����TYu���~8:��:����G(A��!о����?��\�F�4�:�
���e�`��7��4��y�W#��O��k ���Es���Sp�y|�� �*!j���;�J�Q�ٸy#�^�!M�:@�21����u�dķ̉���J��JՖ3�Z9i������I���M`e�^ޖ��lj�?�s������wM։3 [*r^�5VAR�hx�V��1�0�!��6���/���;�]�L1��{���O՜J�g���[<@O�D��HC�zz3�r��r~��a���,���zQrN�+؄Ĭ��x����)x���4B���A�v�3��`VS����jK9����?��C���w��ߜ�,����X���tG��WZ�n��<� �؊1M�&�2_0�ܜY�F)����C��ri�!O�0�\��c��#�v;t)���eIE��L=���:���2KKbl�C���R���z#p(�P\C�������[d鋤(j�6�f[��9E[�o�1��o��k͘o��Pq�����8�;�X�$��ӆ� �����U]q�;L�빕/"�%s�K}�9�ky�2���k ��^�;��!�����=L���� B��9GDO_��j�B�.`	�ҁRA��d#h��yx��%n�r�鄠K�Ip6t�R��B0TVA��pP�|���(|z�ԡ�݊y��ԄFEX���_R.�Z���;���������H������ճ�!��?B�ϯ�������yN�BĘR|+��mL������H`��z5v	A-�4�����xb9�q�p?ի�\��B7�"��rL�'x�8!7���4s���k���S2�]8$LDW�_y�Tض���R�F%\�nf�8�(�n��ݠ��yT_�+;�ni�kQ������|�OK��Lu>*�l�mu�f�u�|��qyO�'�Gh }���J٫�7�����~O'/Ĩ#�^JJp7�:���jy�ҷׇɿP��=�E��e�'�ߋA�����WQ{�K�1j�Dু�"AA�GQt��E:xm%�UT�!��r�wO��,y,�6�V�K���y����̾��2�pb�#�V� 9~p��oŰ�G��aL�좿�"�{�]�0~�턓v;�xb�����ω�1�@�Dc�#G���e����.x�Ѱ��#��xj�s����/	4��8G��z��:rEbSI1=�EV8_�^�Z���[:���\�"��T]�r�0+��ZmZa��p����Q�_�<��H��1b)�����$����7�V�_T�g�R��hjZ_�6ԙ(|1�������Q��|��6��fv��_*��{�-����� ��͠�)�jX�6c��e5m�(�4���f��@�ᚼn��X��r�%AC��*R���p�c6�ف,�ǲL���m�&����y'�;��b���.�oR����J��WD�Lr��]A�4n��<G#3�*��d�[ٌl�r�މ�^ط��r��T#����0�P��=XJ�0sz�-l��'��9H�g�}}cC�+I�Z�� �F���Z��8W�}[-"��M�%�����m��p��R �w����n>"��w��64:��6�� �ۡM|����	�L�Z��s��^N��xF��@�d�C�.a'��@Tˌ�ֈ����-�p�"�8��N}��kN�ӂ�K��c�7)K']"zz���
yIq�h#��rD�:2�-�GlG�E���hɰ�vl��]-�E."��t��M(.Q%HD���m�����~��?��S���N������m�ZcZbܟ�3�9 ��N���x�j��W�[}Et���]	���s)�_�d���7�m�m��|�V1x������M��eu���c�*$J��XP������.�a}�󫕪ɭ���9Ix�G��or��� ���MK�!K������:�c��pF�P��f%k0�F'��V�0Y���=A��E�8u��[�_�X�j���ձ���f�1�8Ȇ7�'� (g����4�;챹%�]4�����j�v��:��Ph��hG�l�k��9���\���QQJE�ޢ�I?�R�1h�C�8��{��a1�Z0}�X�bT�b>�R��,T��\���>~I�*�FqU�x�g����{����Y�a���"���и^1�X��p|
�b��'kџ���-��}Շ��"뿗M|G�  x	������)";}���Кj��պ�������n�`c/�\�t�4fF�;���u���������]�a{�<0��? ���Re��@�49�/��R�a.X��.��5��[������'��~ɣ��"-vT���i$��%�I���_��/s9�7%���_c"�����_z�E��(���xAa���H!��p����;�C[8�-������OgTw]X⁼m�]�|���P�
)�4X��.�X���$���zP=rz<$��d0qT�缱�d�.�������z˖+u��~��׃�6���� :��R�2<j5�o�7f��B�f��j����ݺ��'�UA���54���R���yZ���k�ӧ�>L���p3G�>bŸ�#_���$I�:���I��1��f�*�d�{`�=��r�$.�F����Uc�d)��0������H�p�Cf]j��l3d�ҙ������Fvf��;������tr;#�e�h��j	y��QP�Г��*�n�E7���z6#�(YHZL_�e~nw��@��A��0H�5�*��s'l�8k,_$��,���Wڛ��vE;���b=Kn
��,籚�E�����׮��w���ğ��cJ�������=���י�}��a���c��TF��p��[L�6��۞+��e!�R��po���P-+��u*['+�-�T�k4͚��oy���Ty�J�f�T	�`2.{�j�`�LFӷW�� +�jػ����Z�=D@��Q"�.�,���%v]��[��*ט�N}*L�o�=�K�FX~Ey��7�1Ż�&Tя�v6M