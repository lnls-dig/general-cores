XlxV64EB    455a     fb0"�}����L�le����k��	
4��A	fTCFa�uЈ�z�JwV���n�JE#��{EHv�$VAI�܄S�"��]p���+�$:vԴ�Dcop��]�^��@�_d4��v�*Wl������L�		:R�C�;+q�r�;"gGe"[i̏Y@�3�K��z7�
h�'<�`�������ʓp�j��)��{Q�����Tn��+�	�DR����h�v�������z���q����Y�5 2P�������"*H�<R��`�T�"dEC}D�D�%�gWG�}{{�ș��?�!����5��֝u�@OQ�(��|�u�C���*֠"�5Ū��A]i�_��)f�L��Ͻ���j���<V����J��B��}������>�}���}�ˠ��-o��C�sq;1�^sا� �n�0\+��.pˀ�a��_�>�N���a��~?%�ζe��F�L4�TT��6�p�Wk�4�����.e\n����Pz'�xץ�dT�N���7)��ي˧:�E~���)�?�?�	�-�WFCLZB.<R�q4�ư�k��D������uZU&ȩ&�:�­���8iG�n!���X����u�4o�]r&�h���$8��_a�/�V��B��������#\�U��[,Q.IUPTzQ��0�9s$�^Qoӂ0K�W_�-�tHh�#��rx�v�]\[� ��Yv��HЀ��Ƀ.�7[���?8̴#����#��p�FPݵ�M�!�>���k4?M�w$a����1g��v�,,��qcn
d�˰P�+��!f�#z������O�$.�!;�U�>yf{y��Z��������uXT)��tì�+��>��Ȋ%��Xj�T��z�;3 ��щ�-���׬}��&�ht�:2o���K�h����z�Y�݌�
���Eʐ�P��N��߷�I�Bv[�"'V,�E���>��h`զػk�P���k���W3��T�^���H,����^������e�n��o=���<�Q�ጉ�2Wi�ؿa�0�l'�\��zL���xnD�)d$�����x�:=�=Km���\�ԉ�^�.i�^߼�����YE���opJ�g�j��M����sD[�UMs�U�!mxj�~�Qf�g��E�m��9g�S��k-1�r��/�Y��z���g���93F���յ�Q�0]�R/Mg�������GY��r�Լ�?d�0fe��E4���5"��^��ke�%s�	���K-�7�p$d2�v�nL�a�`�i�梑g�|7�Y�0x���(%�T9�u�s���9�S�ز�����EQ{����!-�N�+:b=�8�D%�B?�J�8���[�;>�w��>�>R1�f	Nm�[������MCm3�{YI��?\�n<����UD��I�7)�L6�ly(��Pk�l��m�����˚�aɺ��ؠ��-�=l�+��7�qt�tH�x�
%��}`���ۼ�8��k&�e�7L�����6��A�b@����ݠ W�})���;k���5�Z���{��������@��Q�M킖��+��}a)��2ٲ��P��¬�t���8!�]��,�1"ŵe����ۤ�����W�P�&�L�����<0@=
/�o�F����!�t����r�v?1k(#Lp�p:�f��^�u櫬� �k�
q�~�
1�
{1n�5l�j���&���,(?���ђM��錃��\�]?*_�z
�؇����z5�$7�>S�Z��� �,1���J����^#���$(�-���h���M;����aa^���٨���*�b*�Yy����溺�䨫��E̸�j"(GŎ��^.�H��hgБ����ks�^��	�ٲ-_N=S뎺/� v*�8X��&��};�%��l$�l�Y~��i�U����3� ���ko�d����ʔIL�ۈ��
v�#�E�|��
��;�^��G"7�!gz�i�v�o�^���{Ĉ��T�HB�\P�U������,�+�����!�i4��(�/Q8���Ym����y䋅Q9�]	T�Y�HA����� �i94��?ҕӘ9�H殮�㫽q(#�K)�U�^��;��^A�٪2g����ǀL����Y��gp�:�Ʊ��L4������'R=
G'`���\�3%�]G�Bެ�4�NM7{�*�_bF���y�f4>�Y��Yc���A��D���Lb����)��O�C6-����h	��:]hO�c���K]�v}�%a�iT�p;��ϨB����lJ>y�H~�6�J-��p�����e�m��Ԉ)���H3�L�(j�G��X �0�n�I1إ���yȂ���s�aIC�B��>���·i�"� e�������9����ҕ4�?�6�"�=�Y�Mu���-�zgW���p�|��)���)�\s��4;�k."����Z������bR�6��]�����.V�Q,*�E���'�z�S�%v(�F�8_zV��,��� 3瀏�_��ʡ���eyZ����Q���M!�9�K��3R�XzD�W���[�҂1����N�|���K�ß�S��(�f-j�ط%��n�R͒#��*r��S�3{U�ܶ���Ԟ�&��7J/�Įk��c��/P�;I�f3d��m��o��`T�;+��Y�M\@s�7ddn�H����٪�]��Ժ��;`jo,�3����C(�Y�)����˪&|�7��ѫ��
��	f�AC.6�Įs콃�;�e�M��?����Ts�[�@}�����E�ZZX5ݗ�}��P����7N��?ؼ	�:F���~�A&�C�O�ש�Xl��eI�~7�v�~L@ת���ѰQՊ�6�O���e��կ^`�¾cfz��H��9r�Sq`9{'����W�F��z�I8V��0��n����b�v����+?�x�S��*�66�#������$��~'1 d�]e����v�NU�N�
�gW�|ԏ��k���a���B�YKH=�}�Ҙr�?4����/]0?d3�4��5	>�����s���%��E�lD�c9{���  !{4�J� 1N��-�	��Ă���r,���i��S���K�,Z��H#��P��ؑ{��6E�z�s�q���� a*B7��>�D���Z�����JᐦPw�%�H�k�T`�N!��ʛ#;����n�X�B�Q-�1�\$���BLz�kDŻ�ցt�ʘ���)�{�Z���s}���.�^A�NV�[p�����_�0[�<�����%Sk�Ԕf�+4U��(�[tr	���Q<�ё�WMś�zt��?>��YZ!�|{�&I�윳��}"�e�o�jx8��k{w����x/�ht8��6Y�6�c���W���ST��4f8;ϰR�n`F����=@p�p�	��Mƾрr��������H�j*��O,LV�`�Ƙ���,s��a��hc��/��>7��@�i9��A- �b��3�$i�!��p�}_VrD"̌�r�Ua*����AxFh����]C�z���m�h<WM�^H��!��d��*��#Vw+s"2j����͡��c.�f�����=�J�-��\�;�5U=,��,D�NO���n8C��h�焒h>E�O�=)��á�4b��_Uk�J���<���_�/�(�����$~�O7@܆ɓ�x��C��oכ'f�âV#,Z��|"�w��n߂DW`�D��@������z��l�2_="�IҾ�ė� �U�
;�7zGK]TD�Np�v0�y�����O�Sק������1�՞�+�p����Xܼ�0�In�����i��P� ���+��~X��gky,��<�JgO�|�mX��d%{f�*4������������}+�pb��h.�.+U��A
�F��&�2��o�%�:�Jֈ�{���m�	