XlxV64EB    2ebf     cf0�`�V3��|���Q0h���?8>\0d!c@�V"�K�Z�%���h�����a���w#C� >�Ȼ754R�N����^J��Q�:t#���$B��C����2���kWR�2�<�����q���ϞH�si�7#�D�L�yA̛@�J�
��x�Z�4���G=:%�=�W�G�i8���X��{E���{��I��
�ނ�kq/��ٽ�������򮙖����	� f7?؊2�f�#,3eR����1���霷u������?^Q��:��!�d��`��>(4��'�$4N>�pҚ����2�<����5�_rMmZm���li�j9���v(�6Ĺ���1 �?��!3H�����V�aB���ʁ�[��Hl�{����U�L��N4١.ˬ6�I����8B,��e �-0Oe���a� ɋ>k2T��ٶ�<-�prr���"I`O]p�Z�����k�i?v�3���(,���P�y�:f��f_&�_�~��hM�D"��`��=�/3v��V�rb�3+~���D�jV�� D�5��e�A��1���f{'K��&\�Ӛܭ�Y����yTg5�R<4��n�M+r�!�ˀ�T7���l�a�����䬜b���>L��FY�a翓H�i���WKWu%�H���O?����
�D�}#D�~-���.�m{�cّ���|�4�T�����&u1����P>��r��.�.k���%�t����2<��v��F���z�VE�Pa}83�-����=�{\����;���c�fKsT��џ�AL�2��3��A[7��ü�~�j�.��d�D2�*�!��dN+1lq��@%S]85�o����p�U��5i�Ђ�H<�c��H8�A���dR7F߼1�8�������s�A�!�B��C'�a4�c&B%�L�&��������. ����=�_V�B-�O|�J_e����ỉ[��r��Dj�W'8!���H�Uiehc�,�:�3�Fo�W���b�>�1~ǡ�h��o���j�p��
̔���جJ�c�i�D�_��m��zzl^�g�8:�Ɨ�E,f�|����-U�FC� ��@*rȢ�2<�2�����ؐ��t�~���@����,�Q��-n�:�����ߟ�Ů}	��t����x��x�>����� ;i��UBT)5��~gF$�B��pof�	�j�6֍r�A��\y�@|�q��o"����3��f�*䭫�'�����t������O�'
�.�6;\��ZHM �@�t�<߳���`;�>����K�@��v��l<�� �����D�R]�!���aXY�̃��ѕ#Up��\�'gg�ǻ떪��^Jg�>1��H���gq�:|TsѥU!�]�ڎ�.��B��eU�ޅ�E4�uTJ��� {�qL��AK?C\��L��驤ӳ���q�Y�ٜ��~8y;�h�J��}��K�G� �@]�L���&#a�T�}w��O:My��_��q��7�w��oD@�.����U;z �s�w/���0� u� ��ʗP+�1�������Qp��p��廃�>������EF� ��˯��gŽ�U�����W�����̻�����U.P@t�{K�1ێ��o�������,�W�k]�2p���{B�j�G���֬��.�M�{�_��x�E���r�L�iq
)$��Ѐ}7.�"�;�n|H��⭯�^�?FU�±m@��Y��|&���3���ٷc
�"?ɴ��bJ�Ij5�K�>��\R��&�h�9�K���$@�@�l�!�'�1'sډ�CW0a�(�Z4��M_�S ��E�!�Cg ��8���M丞S�{���������tx�������������!�~C�˞��U"G����K�]`gd������j�9Y+��=���d������B/��&�pت���oD������B��������9����� ��p� ��`����PGPe~��{_���58t�/��f3u�o���b�󀑹��O������
�8��]��t;#���YͧN-i�<~dO�V/b�G���h���y�u���k/g?��	OZ����
,{�� e�^�2�jΧߡ���P���z��+�m{fU-�61�#!#��ܪ,ɲCf��9{���z��e��7�����@<>5� ��^(k���������a_�cMZ�=y-�u}%��y�x�u������L��ۃ��5iW��Pk(���BCۤ|�M�	�"��AB�@po���D�؜��\_��3�/�@Y"�v��da�<O�����]�'T��/�"�-̉����->��;�0HE��8l��y�w<�R'�K���������MϾ�^OS}R���/R%���tCH�����XG9:5��V��/�F�Y5�a��Y�,�Ze
.�hn�ӳ���B9�Igw���r8���ŏ�� y��n�" �R���3��9�����n=���j�Ω$/��pP��V������ �į�+�g��[{����Q:�h`z��#�f$���?�"	��tv6҃�h?�A�/lY*��s��R�+��x���s|�p�j�
JIB˪�7����b�c�nӐ8���=B��KCA#���^.q�����\����{K_��O���e@=ߦR���M�z�k
��`�l'��;��u>Z�.g考�ʆ��g�)3��x��̆te��� d���7,�@��m��5֢�ǣM������EF�_����t���n�ܞ�Kb�����;�>P�QH���[����!��D"@U�iD/3�ܺ#��l`��j��q������UU:c�p�;���9/x&�=�}c��0���^[VN!�3�
�O�
^�|�xL�ⶋ��fR��� /��y�iﻓ�.뀿�������I�	1���� ���&�K���b� ~�9TI�>��j
��LɌ�w|$5�(������U�D�R��%����S�mxm��Rf-����Y��ը���l�vUkQYQ�mk��1^pB�����C�S��0��C��
tZ.�ן��_{�6���0���e/X{�o�	�1mS��l'�d���^�L�=�9��M�?Z 9jcw�g���O�Έ�PON�np/5FL�!�9G&�iү��0��_Ya�@���˓r�fG��/�\._�@�&yM$������ӡ�ηC�8(Wb�J-1�`YW4�(����