XlxV64EB    fa00    2030�p��n�@(U�	q8�IN��J��56��7��	"3,Nͳ\�P(ށ'vx���NⱚT��i+Pr*�./W������?������^����8k�) N��[3aW�~0q���u�P-^�`M��!���U�	15��ť(�%y�s�+s�g��uړo�b60�8\�llk��jD�[@v��e��$��Yŭ��I�/�B@mg��_0�)��Hg�/�~�-�MUNwc��X��)H.�ᆰ?��Z�y�!�!'�b�(A��a~F<��� �?�~�Jv�|[9����.�z22,u�1&&̦C3n����k����[i�;@T�4Aj+��Mε�|�w���L�zn��x�N&O�D2�?�<�/�9�&��{��+��KS���d3rrzc\����q��1���&�G����a�e���D���(���A@�h� �\$�k�3~���k���{�dȏ�~�p�̰��+��
y�{�a��PG7� ���V-h�.��� �@;[����K�'����<q�WG��$U�t�;�$`�\�TAZ����Ef�X8�L	�9/�*p�TgS�f��Y�媶���U����<�b�d8&�Io;�����y�w��jkV�"D�O'���]/<)��̧k^W��
��j��2M5`�dxO��r����J��#}�1��������i���΋�2Ԣ���1��5$<��U��L<OP��������v�n%5"�i�9!�C��,�"ٺ�G��}.�E"�c�9*�J�^��oNɌ��Fe��1�ǀ�z��!�ݡ�!�?`L�N�X�|�3�	���ˑ�2xt�F.��j��&��HL�΄�H8¼�,Ş֮�郶.�C�*ըof	ff�ïm���3!���Zb�+j!������0ֲ�h��6��}wS[.��|�>_u���P��/~����d6@ۻ��\NI�0���� S�2p:��!�t�P!���O��c#c�a.S:��$b��.�Y�������RD��H=����!��^��>�(��͡L yMf��p� ==,kC�W㩣c�ǟ�a�O^�r��𾵰�Q�?��b|�@%d-���}
�ٸo ������#�� ұ=��Up|]�2�LU�
�9Y�h�0v��1�75���d`<_���y��H�9��@$�J,̟���I?AF�F.�8!uXf� s��%����ACK�٣3�	^3��.��Ƨ����f(��Y7\���gc�Ϩ�7��8�K^�����p�<L'ΰ��-/��2<����˕+���*�?����bX�����p�u�����j��?4�>�dY(�-<��a�X�2c�)��Dߧ@G�r��v�F$�m�hӯ�L�$���� ~��iRK���˴kmաg��(dYe�y�6�;-`g�t&|�b4b/D0��k�-��ϗ��D�KL��5}��bbp[�.6�=5﵌�O/Jd/Ks,/ɌiY�Q����m������!D��Ϳ+Z���c#���P��,���.�i3�DI^Xg��å�K���8���B�4^*��&s2�3
��3�m�r*��'/�3��d~>0J�)����0E,��
�Nտ0kN �eQ�!-���47�_f.���j&m�Μ�(h��Ya��V�N�a?D	-]PBR�ƴ�c��s˺5J�2E�O�h���
��t�d`y*5��@��j ]�"��oLȴ��u�>��� �8�<ᆏ��-&0�@r�x��83��YĖV��R�N�����_w��S&>�%��l�x\}�4L>��sC�M��KF�=��ҭ�(>k8�xb�۠��^��,�T�#�-&Td`w(����;t�9�Y�ރ��<����D����t�����mUy���M��*h�GM+n�4Q9_���Z�+�T�Y���b4R��,�2�[��s�qii~�b��	DOq�+A��ޜA���@"�L'��z�$�sR��<��uUb�t;°%�A�o{���ZBЦ����8�Bf�5�t��8���")�=�-VfU������z�U;���pf�~���&2%�W��TRhKd�[݆���LT�����1T�0;��}���f;�X�v��%�>?z���i!�L�I7�C��$,k����+�qm�UD#J\����E���"<}8��I,���qh3��޹o�ĚF�E��cKԎ.Li3�'{a,��r��#<R�k>��`��r]��"b�H�*w�k^r�^��m�~נ�T l޽���
���g]���#�{Hc��� ~��9ɔ���W7/�>.��nq�]�J�m��!�k���'��Y
��7��r\G�/k��M'kB}�� %������Ӊ����JPq�ݞ���J $����bu*^��^������;���O�k�?�Ђl��&�.a7�>��䎇����Z�!�v��6�<P�Ёn����D"`�/�#�h�_bӥ���F��-ox?�M�l<��/�n"E����&�� �?>�0dn�wÞ��b� �f�ܵ�_�@3:���l����7pL�s��~���s8#�ŷ G��3�͢"� Y%�g�1�2��dV����_�j>W�|���f>��ge��"�-ę�:i�m�W)ӡT�z���/��I�y�����6'�G�]0߳�1���NBBRϮpt�I�� {/~{DX1c�'u�š� V��vj��������i����x%������|4�`y���)��%�����6�J���O��j�g=\��+��a
2����<����O�{{\��hƌ:��jE�Uv�?J��z=�,9�~}w��v{(�� �D������ʋ�1uMZ��vd;Z�dM�-��^�F�e��'n�|�ρ���u��qt�A)�;s�h��E?�9��7�K�ӑx���Eů��<7�e�la�zq6?-װ���c�ũW��֐�1N����Cק-���&���!39�OH@�A��r��+�m޳��"Jd����8����{��WR�S��(
j��)/��;7lAy̭�-��*`��o�y:\��1i4��J`��l�����5V�gu5�7�n,�ÝC���d����z��
�-%�p���[��"_{��.���.z?���-7�b�x��Tw�;�Z�=ɯ�2�ϣq]0Q@�4�Cj��@�S�}�	+�$�#�]K.L�~�ǇR�e	�..���j�zzױ��x�ogV����u�R�v^C�1Q��2��O����/�5M|�*l<�F�7��f���3��84�Bَb�	�\+��+Ѯ[��1S�C�Dv������N�*��d�
|'�0Q�+χ���z`]I�T�jY����a��	@�ܗ�,�́WB���.�l\��]EԍGԠ�i�꧊c� ���M�ZAN]2+U\��q."�s9F�̠2h�+�T�BMS7?^�F����oz�9�g���nK��F������%
�����uDvL�$��7�JͲ�ٟ�]��t���ң;���nutؼ7���o����9��+h��Q*�aZ��ܹJVP�"r�����Gc.�6�_
�F�Y��cվ���A�"�nh E-����O��-s�4 �[��e^�#+��.��N'�]��[�"!";��>�qa3���L����E���Lk~3c�Q��g\r���уS��iI~:�\	�^0���N�-*>�����J9�.��[1��˱�E�/�����A�����S a�����^)���-�N!�T����=�vv�X�9�Ə:�8�Pj�hu���$7βh#��o44ۏ'�5͚̊Y�}�b�S
NSݽs���ɢ�0�����qd��J���
B�K���t���?����N4�e���F})f�=���#���/1K��>w``R��"���#�d.�"�a�%1�G�|�����\����JR�@�r% 8	�Z\���n=�0��N�9 T��JY�6���|�:���142I�*�k[�:�]� �^GB9��Flis�=>����Ks$ɜs�ir��1/wqjz}��p|[���Nz �k���<?�@˘��NG��G��B\�|�=��x�5M��?�i�ćJtaISA7���d0�-|�IE,(�4= ���_wQ���ı��	yT��Y/M�a/��m���5����'CF��g�*'�ǞF[��sG�ԣ.�$�����;�~1���n]����
�uR�� �6�ė�]�Z�N����X���Z��"#��Mg�n˞^0�S۽�!%�4��{�j<�~�,)���k�)�8eLgrvߊ�7!W�9$��-
�S]��P�`1ظ�}��K��"�u:�6Gz~+��ti$&�GC�N ��Ҁ�����r �f%�7t�0}��8�S0�z����B�F|C�G3:�*�g���8�F��2�!]���y���4�Ӿ��)��H�Rt!�ncp�F!�N(�,a�1� �\t'|9�Ʃ�:�S�����gë)3���d�Y�0�Q������N].Š�KB�n��R��_S�j.�t�#$���d\U����މ�#	��y��Ж�?)0�vyIN9朓�Qg��I�|�(�=�c�����#����z<�pPM����vB
��}Ri������|�<B�j=����0��UܜW���zY��ѧ���'S�Y��~���w3���\U�|udR6�[҈y�/EL�׬�p���<#2+�y�+33��J?;4��j�	d�ֵ.g�A|��[5��P����V�VpWU-cρ;��w>239��ś��XT������{還���x@�|k��s�fh
k��:G�J�X��h�l�۪Z�J����H��$���d�n�g���Uzq=Z3�dyB�p�z�X
/��B;q�`[B	_�_%\��K��uO5A�m����7
���ߚ�G̗�{�t�YU<�_I�a��Jc���E3*�|��퀹����V�.`�xYG>C�]�h�I �����Ҡ97e�HT	�z��T2���\�8/�Y7����2J�Ȝ+���g���|�h��ISG����j2|v�5�V��)�'�ԱK҈*�>�����u���b���J��h�9�ļ�M�i����!�L���2���y5�Ɩ�?"%�]�^.�%6rPp]<�3u�� e�� $[�A�~
��������;R)ϡ��hd�k#?=�w�����ź1sŮ.�M�����vgM�ˊw�f����s�HKk9��=W`{~�X(��҄+��sl�i��3��U��� ����M�i|V��{�ۏUD������>��4FA$r
3�*�avc�泼�b7���vN�1���Ȃ�*�7]����1���8z������p3���c
�j��w�����ȁ���h��;ъÙM o�'�Oi"gL��lX&�	�h�>��4�ڡiyWe�S� �Քn�Go�o�=R�YYr67���>X�&z�P���<�c]��S�r�ifM�q�i�(�BF�q���7�t4:�>���Xu�QAc3��u���R��{ki�gK�Y2���׀ʣ��������`�F&u9jԊ��,H���#Z�P�&Կ[s4�K�����t[�c�5������/���V�*uV`�� ���CG��	K���)���4{V:*s���1GP<xʈ�1���[zv���:�Q���.�=��0U�~�Jn�#��Zb���.釹N�Zԟu��Gp�xi�C%X�P��{�!���8���i1��Y	�}>
���	�g�k5hen���𶍣���M�3�H��v�¹A��x(ȏ>���9\�`I}��j��6B�{ͯ�"��-V�Jݰi�|�k��$axi����$ʪ��M�x�G6�(4��|i@�7@��y�jf���,Z(5���Y����k�_�H�L��WF�s��M�tca��(G>�A�6Pg��a��R���쬟>���ٕ����~Dt�ќ;?�%9��\)���Ո�C8�6�0>\��(���J����Ky� N+�N����}-2���P�q�Nvt��z�p$�'$n�hD�F��oJ`�u͔�:s,��TfW.��'�0Z�м'�gɮNpW�S��n�4T��c!�W�/v���6G�"ς׽�yf;pX�d��>|�V�X�C��j�TM���.U�*�6S=2H{5��D
�J�J�����kd�߫g�����!��5�Vc7��g�5��ϝٟ*
I4�� �Uo�D�[�7�ago�0Ajr�x�����=O�Th*�������Ƈ¢~!����o��]�=��rw�y��B����p��H�t�#�+i�Z�ϟ֧t��\�41V�6��>G.����ė,)�&�E�(����T��;w9.�����vz�<��`Z�����-�A��`5�$;m�����P�Y}�zC��e�ڌY$�_%A�#�����8�5�UD1�Z��n���������Z�A��YxY<�*R@�#�
{^�ot�Dɕ���l�]�ÿ�@U�k�2����]&��x0�*N ���Lv1l�P_�3��j�熫{b��-ɘ�7��CW�i����,CE�4:3�)�5�[ܯ�Q*Z�����&4������"օ��u���,�����\d�	�1�K��p�}N
!S����*2�2B1+W�|�����H�$ԅ����ɖ�W�)h�I�� G(ik�,~T�eW���$�?��S?T^�^�*����,�b]Tkɚ'�B��8B: 8^����Z�Zeہt!o�mi��C��3��@�`��]��>fN��?�Q�x���ޗ�����&����4j�eH�Jӡ!Xu��4�t�"�UM�*.��M�]Yq|���[�G.���p�:{6�(�D���5^���~���U ��pˀ�>R��w�0�c�,��s8��+��#�oSG�bj�r���@V�@���ۢ�"�Q�<���P �R�ֹe;n銤@D<#
����l~J��hӑ�ll�>�bW����=KM��D@�߷�T��7�5���ۢ�v�ѹx��!8W�H�R��7Tp�f�)��~�ςn�`Y��i@g���+�ar|��k2݂%$�;��0I#����P��HJP���݅V�(\M���}�*d&�F$�R���F/�6���1fB66��MUs�!=Y@c��V"�v"#�q�����H����J��p�7X���ן�|ͨ�C�s�#>~'���SY�JiW *�i���n�J�����X<�L8.tl�f6�a��D7��Q�2�ϋ<�� qI�X�# _��'�ST���k-�����rD�!K�vr��ȍ�H�I�4w2t�Z�!�}���OO�|jJN&lN��~�D�Z�ad;�W&ڪ�j�ϓS��������4FK����X�$�{�;
X+l����������ejG��q$��	-�9��Wd��o1��n�DRV?0�}�&�1�J
u8��R㏽�ʞ�CЇ��	z�C-}]CQ��'@X������^=�Ŭ4my}�9����"Fز�t�|vq^#�X�w� ��^;+�~֨��>aJ�۞��7O<�&�����@Ts�L�{HekV(� �5&f�y�-k
a�D���[��/��y��OR&�p�wV�0X��{���e���g�@:�6�i�]ɖ�S1�mO!{��d#T�D��	��'=�8�/J���*y#����sJ֩����a�ڈ�	�#���gsO�������K_8%�q��r~DK��V�oD��;���%�Sk�U�ͅ��,/��vw�X�S�S����a�v��ђ�Ee���	Će�ܚ�eߴϘ�"�&��SG����Xw�a4\�,��ErR���Bnpd�U%n�d:����kf�� TH��P�
�L�9Q�[��� K�����	��������u���P9�s����F
(�iF��S0��9�}�-����y3�jrS�H���h
+U~�����"�`����c	W�j7�0Mo���K����(�Ό�����C2É�K[���hV0 뜁�1��v:Z�<�O�|�XlxV64EB    9b47     ed0�
�d#���$�Z��e��^J�$�'MS���+^��%���MJ9�D���� �t��ܖ��p9$qdt�^��\2A���ѦY�`�:*c��0�[TP��û]��c�l��,(8�:��5H�ɽj�yV����T吓���g5�y��XD ���<����/����+�+]����+�2&q2�"�9OڥҪ���(���%~�z��%�&�ìE͜qmU���9�l��6kT�8e�B�,�B�ɠR�&n��" ]S�tV�`�HK� ���Np������,k�T��9��W���bwx^�Fi�@		�ϰ����4���������fC�p���[0P(F+�{�2ӪW���}R)(��B���޻�'N�j�l:���EA6?0���t�he	̦� V=8(��7��6SA��rV:jD�+0���7 
]� �a���u�Z�gw�g��������!.�����ZЩE�&|�����I~}��%��\� ��y�F@a�e�:6خ��r����������$�N	U�*H�p�Ir�+�~+�ς�#3
2q>�@���3��o������~݈lO�	4�;;'7v��@�όT���U�U�¯�:ȇrO��Wε��u�h4޿��O��1�JH+n��Q��FԚyK�i��)�U�H�(?� ��ܬ�ȿ󗄁uP�$�TO�·���f�7�V!H*��MW|HB��ȣ��<2O8��ﱌ�V�f��2G�[b�{Wз��^�<s\��DeE�sE@����^�G�����/4�������$"�%�s�ԣnɵ˔Sp��#�Y�DW��Mx�d�*	b�7�Hv�����M8�����&5��(?����~Bx��L�Xr���V��(���O�Ց��jr��3��Z2���jD�c3����S�n+�Ż$�:�)�DMOg<��F|��e����+��K���4� a�TD'��l2r����Uړ�B���9�N*
4C��~^�ax�ݏ@�z�}��ta�/��!m���O�̻p�Ƴ���� M��; 8�ѳN�>�L{}Hv�b ������פՇ޷�ڈ/RU�Is`�?���W�&9�v�� ͧf�[[<L$t���_������QU�p���Z�rXl ��}|�)��,n��jYE�l�˘\g3?�l�@	t�[����~7����Ax%�����0�mѱ�`X�F֧7@���(M����� I���`)e��$�m/D���&�YBe������~$�G�%J4S �@�ş��É#^3Tp^^	� pt����5���E"��#u�c�4�S�a�'�����Sr�\�X=m�F�Y���1��&-�G�����\
])��~,��v%�d�-.|qq���4�m�^��wʪ�Б�H���~(5���㻎\�L� qf��!xF������W������鼩�"uIр�U�{�c����J;�W}�E�y1YV ���J{���?�
�/�3����޽v�+��L��������W.<H�Bz:�<�w�2g墡�%��f�L�İj�q��Id��>��#A�,��-$�³�am,jS��\B�6$g�x�y��70�D�^�xܙy+0�5�5� @C6���#IPWM��srNh\�?���E����b���#E<���x��$^�yX}z�{�=�ב��i�R�W�"�*y)�楸H����at:Mm�#Q��TQ�}�}��W����.��J�9�4����P�.�~���Jf�!8Gl`���5�*���s�EE��"��\�Bt��[�_���b�ɮ����~��s��î����vT��		�Q `���B(F$.��܃���0�=�o`�vc���Q�7A�w	�����_�Ֆ��8XRx�k������e����-HH��~֢ne�1�lv�'���5ᣨ��� %����&�����C��wu:	�nB���ga�\��{��M=�tڠ7����fy���IK���e��=�u1cߐa��2H����Z4�y/�.M�-o*�I��Fm�XYbNm�@����g�&����T���M!�]؝nn�a\3�Ӌu�Y0=u.g��VC�;��.7VL�{�g:�Ԑ��6�]^F%`�Q' @J���I������)�2�ش^��aVe�v��F��x>N�*@�v#�X���d��\o�3 �vkZ���z�rD�{nZ�6v��w��S �)k��vٛ�g�x�n�zްʫp��}��3^�~N����G��4��\E��S��݉<$�R��X(�h�νD��%�hI�G)�������ё$1�lq�b5pR�6Ex�#���C�ɣ�5N�Q�d�Ssk4Y`�Vo�t��	ja �p%K���{?���[���l�CVz�<��£����2~�m�P9�؋3O72��>Yx�����`8�}�2D>B�V�+��W�'g(�A��[��4T0���o:O|��*��&Dr��A���7C���[�j�R�!�&=�i�x��3��?�D�%���&S@�uu� 8s�׷dΈ��sЭn��~��G���|ֻ�[bu�c+��r��@ҵ���l�{&�H��bB�⢄��z۹N�%0���	a˔��xM��rw�j�:y��L��3�?{V����	S-�E�8R����QF��ɷ>�,4tk�����;X����?rxp}�C)ދb!%���w�Jt5oP�"H/����<K6�|�mQ�����[bd�`%�Z?"	�n�~հ�R��̥l��˶u݄��R�w���S��T�P8�w�v^�k
W������.�0βsߘ�VS'8X���BC��1'�PQ�<c;ҙnv��^�~ۨ�#Lr)��j4�Ik���`��p���B���qK?�JY�Ű�&���e�Ka?��F����45��ܒõ�T�>�"v�̎� �Jt����+���E/*?%❥��L�D�x��UL;�&��#�t���?W�ц���J�����^��j�:6na�X�=Y|�D���:{���a�&&��:�$	�S�D(��R���'L���b�Ť#�M�]�|ƽ`*�a��]H��
Dyݨ���[�ǯ��4�0���[|�$��W\��𹾽��S�s��G����:���y������������:1QYĖZ�-n���Q�Q��i��q���2iNZ��{$�t������*��Lܹʙ�'zK��ձngx!��|	��4��� �WƠd{��p�иլs]B�k�p7���o�G>#��� 7�=�u�s؅��}��M�`�90��&��a�kT�K���4Uh��S4��,F!��Tpv*�b�k� VIui �l�3�$���s»��.�s�y��7��F�	*�2��	�-H`���AB�|k�J�֌<��µn�w�}2�	DN��Tb�̧H� V ;�o�QF�*�J����cA���5�"*��3O20�O &�[����?Ԩr#Z47�!��~�-U��/My�,ȕy�@g�s3+T�Y�s�vS�z�^jse���>��
��r�y5�����'(4?j�)Q[���C�~�d�ld�&)���� ��
��(Z��e��es��3Z1Q��{noKD�\�]�����&'d\",�_G��rsz.׼Ϥk��Z�5�Y�&��9�gO�,���j���`0�B X���lG��]eN�G;H��S��x��2��G��`Bq�����08���"Ǎ޾����{1Z��k���5�ѭ�h�