XlxV64EB    8760    1a70���1b �A6gu��BA�9�DkK�1���''>u#�t"����`ʖ�3 ?md�<�쒫jn��ҟ���4q���է�A�ƍIo4*Q���n�:�
�:�v�_>0~$�X�qc����`hG�U��ֽ�����Ө�vUm��z��zF���R����48�y��Ǩ�l%���Ձ���Y��sDQ������	t�8��pm�����%!�@̱ �K�n�2�:�vvb|��R-�ǋʤS2�1�"3���qe�m�B��d���-E9�Z6�J�,�M��3��#��U��{(_�y&���\�����G=�mY	n�Q]���n���"�ܶ��vGʭ�)�����NI��>� Ù�w�8ij]��ֹ����α�����rua̕o+��R�f���=��\v�,0�S��-��S�oa�Kikk
��=�/K�Vy�t᷷-FD(Y�[؃Y��+��E�!�*˫�r�4�]�U�E�8ū�F7C�S��ŧ���<q��u,B��}��/���ySl��B)�Lp��$�-to�N�D��b���/���^���ńe�YDGK��3�֏ ^�D��I�EtP�6J�N���b��Եy_���J�\;���H.��� �O����F��km���G�	�k%f[_K��	u���sv߷������Zp�t���4C��O�����}O���'��} �Ŕ�:����d7�W�N6dk���Rt�@[��+n�%e��s�k�~ �ƽH���Ep|X[Ԝ��-H��v_�P5�q��vyw���=-�K,�Lys�xr+�;f�6�[̽�~'`&ߑ�r���ZJl��1�b4��v �1��5H��`=�'�i2�N�\X��p�n�-8J���(P����v4�b!���t�KV{5�8خ,5A:*�l����arehr)����Q.�ND�x���7GjeZ��!K���{����YmǺ����J
�;Ov�:���}�'�"��Ҹ`\����?5�����@#�}z�\���u��ID���#S�����e����B�ǜC�7z�}���6�i&>�m�e������Z��h��׹	�4�b&�o�����M)������1�:ۼϗ��d��8`�ؠ�g���o!3r?y���ie`=|��9�X��{S�@G�t0|� ��lZ��K����pu�یݦ��8�,��yP��9Et�7��xϣ�ȯ���h2#�iH��d
��,l�]���m�����BF&GҲӗkZx�oX%�[y�,xx� �"_�,Yz�'���~M�Ϻ]I.�]�́z��S�[�ٸUI�D��76���Cb�s1ᬩ���%Go�@0m���)Ԅ�ȧ�Z�t��c
�[��Q�|~�%��o��ݻ������oŵ��~mT�	Os��;b������Q�Ԃ�����d�����l��3�@�˸=���9֓�tz�%@�1�d�h�5�[��IX*���iw��Hm���R
����U7+��w4v�.W��U��o*8�MF�S�|>1��&a�r+�����!�.���w�ɠ�jAO*dR�{�;�к�hm��vA�3��J��@r{�@F�0�&+�Z��hw�x��Pkx�� n���R�,,��i�tg���� �i�i��KU �Ŝ?�i�n.�5h��U7��1,�zvhe�S
 ��G鶴��6N�f�jh��\��R6�t�!6�e*�9��-�0Nw#�wL!����I{c�����~�I$[qä���0a���2����Jς'��U���`=1����@�$A}!b���ܨ���J$�U@a�;�+��y>��$��8���ˋ�W�m>�%�I�=r'P�J]���~8{�f�k���K2 Z�	|�υ���B����imK�&�z�R��/=H#[��=3��#GqfU	�s��'kU?}�Γ����E��P�\��ǲ�"���Lٕ�/��[Sh���\�+dE��f��O��}�(}����?&]w���Đr��e׆�>�-�YF��4�8�����7!5Y�������P���׍Ĭ̾�j��sr�t-I/�����y�1�U^$HY�׿_�GX�
m��ڭ�9�ׁ�_�U�pdŁ@�t��͝��ş ���pE��b��'R@�VqFz�Y��%�W�5oD{�6�&H����t��@v$�~O�y�Ru)�:{�.=y�yy����f��rb�^��î�zPO���1M��c�U���yA]+C�����:�@� 7j����y���fԹ=���` �&������x�{:e	||������;�ݰ|�.�m�&UA�����ty��"A;!����'����a�� �V�f]6A����$j��7�Y9ڽX�<^��*QEW�6���M���	���FI���k�{��C�ڡ�$�3���qnȎ+ex�<Y��i�u���[��tr}�i
��خב3i�!r����-�E�^_�z�ѿ����2/md
�3{���,y	�\	�Ln��S�Ru�BW5���f�J������{�?(���R�t��m�Rb�X�@y��l��Qmy���\��Ev�k�X�.�E޲����	M���'X�߉�:f[��yj\K�SYx���"=1�t��G�J�/��Vw�=��\��HJ{N�<�����~X��yy���S�,#H��&�LH-�䞫$�����z�3�J`]2l	kẬC�0�.X�g`��.K{e���.�s�d+g	�ZN���	�f�sY�z��2Q�r):�i7�} �pѽ.gj?9�
&��L<f	rt
o٢�}�N=z-i?b^�D�X�H��b�)�~�*�j��(��)�h�+����vсq$K�sd��{�r�"�0��� ��c���də^˃v4P�(t��J����:�6P�3>�ih�}j9��(��^�	B�׷\�� $�h�a�;G,�y���Yrk	��\����D�'�W����(�ۛ�w2c����p9��h*����W�w�J'��<�WϞ����t��D��3s&�����#9�dwW���y��1� x{g�N��N?���F�#=1
�4��t�C�]�JYp�[d�}lP�M6h����tUo��Qm������b�3�Ij�neS�5�Ķ$z��3G�UA{x*��[�̳u�m��Z�S��}�lT���J�$v���%/2�A�pzE$�Z��/��01,O&�[��(h'����1�=j�)n9�wi����>��M���S�ta(6-��;���T�b0�?toP��UEYP�V��*�>4�\W@D�:!��ı9`	��W=�#&T��ةr��.��Mt����l�(��L�Ӭuƙ(��@C����C^�l����.Y^A%�D��zS�S��<R��atRm�b�3K�����V�����c���Ji�J�@�7($�y�{4P�Ru�h�WW�<�0��e��
D����2�a.m)�����b仉��@B� �!&(��_۾��f&�R�������,���+%����T\�N��Vӻ�%�,�t5F+D	���������[�
��D
�gY�R_Kr4F�~�K��<q��n"���]����7V��gvC��M3��w���D2�:���`L�+?�~��2���j]\h(S&�7��/�}S��m�N�3n�/�T��	iST�$P�.6��و�q�2�i>����b!V���l�����U��%���1v��;dʟ�Ŭ`"���L��.u;��\1%��vi����Ɖ�Q�{����>-!�l���_��g�WQV'�d`VLk~n�n<]-���λ���}�L�w6D���dּN����P���*'�X��d�t���Cl�{���5�6��?��S�/j�dj�jd8z�gR ���OAbT%��u�s�h�۴j�k7f����S� r��Ø�;r47�&���b�=��cz.\�<�k("���2��[�*T`dz2�tkpöD�����Dm��"hVZ�[tPD�H�h�ҁ�����=����}�<��.���{��D)� P�<�b/DD��ڭ�E ͅW��Y��<�q���+y�ų{�O��soh��E��Z��Z��2���s-Hj���3n3�[	<��\�/6"���\+UC�sU!�KL��Vf��j�:$�nlnM�o �1����M��l6��~Z%����� � y����n���X�x���k�.��L�ݜ��cQ�+C{�2�^@���EċË�8�;�r	uA���}I�X0�W�װ�+W�$��^3��R�Ǉ���
pa��sŌ�H���G�q��q�� ���� 9��Q(����4)��N]��\�#2�gh����}��\@�&��2]X�N�M"@G�)%w3�ϣR�3�Q��K�M�:��d'D��C��~�s\����c���A�-L��e���c�D, D��d��'o�!*k/D颙Z�p�W���d����)����cg?*S��-4�#�ui�6��Q�PM�������f�4��~ڗ�"!�!�!���=��]_qAC,{�t`���q7�wۯl[��Y�� f�O�t({WN8Hc�w�Y'gr]��bi�lS�~"�Kn��#z��}Z�&�\U�����<�1)n�D��ՃĨB<����%�T�e�Uߋ�pL�lH1��DV6��Ky�1i��Ҝr�K(ـ���9\<��"�Iy���n������sD1�iO���v�A嶴�c�����Bb�G�<j��=�q� ��x���x�*�ʐ�xB�#��c��_�kg���;��bmk�����[i0���uJ���$�=_}��S=R
dB�2���ϣb�;��������c �����v�LJ�se֍�h��!����k}��By�%��Xu-PQ���@��O0_,B�}ZŊ�5O��̃"��ښ�f�Wq��d�z��[U}k��y�8�f[/&�'~&��r�Lk'"+̻������Â�F#3~ǔ�ޤ�-���|��uf/l��m�,]��*�%k�d��fw����������+���^�6�lh��������h7=@q �$��'��-0�`�3�ڊ=�H�xs2OL�+	̫�0��H��n;��hj��S����G7�H�%��{p'�w����2=X�������s�U#�"��YR�Э}/h+U����������ے݀�(���=A��ڪ�&�H	Q꼊K�֥����
oӾ�'7����A#E�����B�bt"r�q�C��{+4�b@�:tn. �����$f(%䧎$E^���&\� ��V��_.N�8���[<tаWC^��n��"D`Wjo� �����C�]v��
[��'�Hki9	�%C<�Gm���㶠��|���(��Y��K�O���U@sx���o��5�}-�`j�f<�� ���x��'�X�1e���ٷ��z�����iQ��.�t���y	�T�9�hb���BF�R�;�
��m�g9�?VHu1��}W�D������tFP]��UP�Ġ͂��+��n[
�)<F�2o��b��`��2e���mH�ZAO�:K��ٵ9`�<R,�Řd�oI���¶��q�_m<�Y�4����ĭaLL��L����5c��LI:8��H`�z���y���T/�DA�y:`x�ӇVF��/�\�|��LMْ;QA6&��Ʉ��^?C���k�I$��s(�q;\¥FI�֪��צ�pC
��"�X�F��w���L~���o��%����]������Kd?{�T$T��7���ޢ�M-������P�ɔ��Yo���|��jT�IU��t����"Y��5o��NRK�y��Zj�y����*�����\�}�6��>w$ؔ@�(g��B���?���A�;y<��:���7�>����i+�.�n�	�Zej����e�NA-T�U��[�EVd��f<���+�T���~�"M�@�Y�XX^�>�����ޞ��#���筰��Ɠ[`�ϑj��Mi�0�^������+2�L�:^3k�02Q���u��u(��澴��)Fl�q����h]TN_] 6������N�GZ�֙��^�U	��]ȗ�Q�����Hۃ�'��:��+�;�1l�A�M�g<����`���oM!C��j��;Jw\S(���uJ�<W��[��W�����(�kY~P�n$��ZHzGհS�}(��v�E�O��x��V�������|2
��6؄+�7rOZl��S���t���q��>y#��!�"���K]�2Y;M:s�s\��{sə!@3����X4V�D������#�a�l�L�4Ѝ6M����L����y;��pf�hKX��E�Z0�~w��~=�Wc�"K�����f	L����e̠Q��~ܥ�B�g��W�c"Z�#^Y�v�+��t��s[�xI�["�w�%���,|�y2��i�y�*������#��2X�Q�z�Ri��\<�{�H9�'���n�m����M��|�t�6��0�%-^���ަ-�r!bWϜn8�o/��T� S�m���K�W��)�x+�d�s�q5����U�#`/L��0��