XlxV64EB    3b47    1040�r�#{��`���Md��a\z��{�\ؑ�ڌ�.�f�5
��@h+E(���� 
�,�Kt2��m��O��{�1	�H`#t�Q͵�����C>�^�5f�b����#`i����eq�� ,� Bĝny;J|�(��6�����M����@h/L`�$��_B�o�B_��(���oH9+�n��t����K�M1����y�J+� �-u
�4�(C�:�L8x�󫺶TJ:����bI ����7L����{�,�c�lJmΓ��Xi�M3�qJ f>2��7���"1PWQ_ݚa3`e���ˬ���lrQ�I��)���56���y_�$�]B
�k���52��0Á��,��/N�Sڈ4�*�w[�����D����������!�3��Ty�h��"�6�ם;wb]���zz�6qG����B��o��dԙl b����Cc�1+n��W@x��<�g�K�E�>w����Zi n8�A��a��~���DoXS�����O]
���m�<���_�t0�.�O�9�bM;
���L�_�t��d�BQ��)=����O����K����s���=�r�KT������xJu��]cB�n��$M[��Zb����������:��y�>9��^"�@��u�Vo�d¾�?��S
Y�G�N��`Qb���<8��;g�O�am��#!V�")��/��2g1𵰜�����)6t���Ù�!�O���%Z�h�BV��Y�<R��� ��^�+j<����62�#U�:N��]����|-��_3C
�����K�pG/��$��%��r7�9��e����'�\�S_hv4�*��o:���8T��l��[�(?H�"�s��W1n`��R$3�ک\{N��^���G�q^A��j�0Ux���*}-`���`v�Ě�p/��b�-���%{�5cD��%e�pX��"J�Rz��%L�.2���j%s�
�h'��&Ӡ�_�C�SBN��8R�]1y�x��2#�٢�V�������u��µ�]�+Pgm��@�H��B�lrE���,S�EL^z&|{_F�����Z7<��L�'f�6�\R@�d�Y�O�����P�-w(歀�6��Ȋ;f�E![��R�B�ጀ{�s����̊�����X��6Y�a }i��j�53�W�X�ZF�R @j���f��c�vG����߯4|������*!}N/m4�����ة��i����lCR6����0��4�鮩�Ej�r�<nJ��rYJ�T6�վ�W�&��2<M
�g�Y�& Y����x`=,�H�b.��P%=i3%�nU�ǟ�A~R�����?P���8��;�D;B0݋v��W[�k�+�ۻCwu}�ZHy|+M���Z&ވ=�$��ϲ\9%��n��P�V6��ɫ� -�AR�c	��\&�6��j���	wj���Q�<^A�M⢖Vu�5��� ˺VI�9���$�#�Sɗ#8}ej��Z�p�549p_3�6��-ý�FQ�"�\`�.U��*r��nc�E��֋f�Q���t�%�h+d�8]w�i��b'�t���͚��w��Y���8+�/��'�|]���6�u�UZ�d
��F�I���g���>��KjQ�d_fڵ�V���Ό�[m�V�J峦2z��F�>���yg�_�%�D��p��rY.#��ۑa��\0��?
��-mם�P?�a=�������Ed�`��}�]��fU��u%�h�'/��%wx��*�8O��%��a�E�����tE���!,�¥q���`F�{A��3S��M?=��V�F|�Pa*zT1�4Xnͻµ_��1���)�X�Ӵ3��K��g��K�Y�_��d.�W�%�_+ˡ�6 mR�"�E�#���y�-�nX��8�dT^��m������G�M�הG�?�ɭ�$\ch�J�:��N_��8b��uٓхO!���$>�B��F��JkH�(O��Ly���CȌF��Y�ىv,�o��a[h��ۧ�?�.3,eSSU�!����u��Ȗ����K��	����qy\m���bA3~�!�hQF��@?��]Jد���!�*�0�W��S��b�7�u�4�S��9�qs�oޚ<k-+lf =����*����r~
�
��y����N������Ҟ_������d�;�F�A-1vP>����E.�]E�}Å��P�`��ūؑ/C���U��r*ka)�+��.�А�9��a�Z� ��Q�x[g�m�]��8��1�%ܛ�v�.}�%�StM�Ih�T�"Ŵ��]�Ŀ����N}�}��M��D�<��-q�5;ݐv%�'r���p4����(��\\n]����4�Ə��b4�&Yz����L��M�ۦ�tx�MB+���q���i�!G E_`3�&�V�,Z_E����e�,��Z���1��d͈>ZC7���?�n�F�1����l)��p�y �<���G9��K�v�.��%��֓��v�{Yf��B�b"���_c9 I�Qp,z�V:5�u��h��I�\�M�o0�h�\1܅��H��W�7�;\�S�8z�AuQ�%�_���
}o��E�Nٓ� ���)��8��.m��£��%����f۲�D������}EJ��f�?�*�@E3�SQ�K{Ӯ `�h;�L�d�FS�Cձ[c
���Zܮ��ެ�i��.��T��{��mI�!����֏K��Qkl�<{o�g����/��yc=s���V,�iB	T(�m��cʌp�Y�������~���ŧ�{���}��3=yq]�����%D.�ӰdS-������MMe��P_Ԏ^���*[m�3��'ׄs��w�iM�D@��
F�-N���q܃s��q�]ZY�S�5w���@Y*��v�x��TJ�4�r�M�^�-�k���e�����ũ#�du�/��������8زa�;���B�_�&-*V��Ʋ�#�{Ԁ�c����z�o�m�j���.�\�T��G,�U��E�|��lhD�/�UYa��%q ��ne��o��Pk�P8�8������Q���{��T�}q�y��#���Ba���<f��K�"�o��Fk`�O�������Y+�9Ǥo.����:38��i��ۢɬ��UO#�l���pL�b�����2W�/3�<2A���uC��]��H��/�{h�d2
�V��e�[�4x��.��l2�fr$��gR҃x���!.��nyz�x�p����md�!i��&�&J�R&��\~{���A�)�F�ιak��O������ �TSя#/��_7AG�$�S5`�,��m��f�A���A�B#d0�%h8��^�cnM�0 ���h^؀���
gG��LAf!l�N�>F�D���E��]/_]�"�`�fh�-ef�~$Gz������<��T(� g߂2d��%��Ϋ�&�����޻�ޗ'��5z&��g�M>
��Xx	 s)w؟��8�GV[22%*F���w�ޔ������:�li����`�S���Mg��o�["�i*sE�^���k���Vk��_3.Z��L�I�9�Y�jTLTuf�.BR0^/��kLS�?�������2�K#��y[�o���(&��߃2�j��"lZ��;��B���'��#`�pC����jǧ�0h���������"������i1�xoWŠn�}$�CVLӺ�ob�m�'�*ܮ�i�Ԯ�� \\T���1 �����Ǜ�����5!�����= o�!3U��#� xy������«)��v4���
��p�@<B��o
�Sy	:��
_�pU���r�O`��k���f�xV��Y�����5�Ɓ�1��+�����`5a _$p,r���)r����1v�#L~+�x�s�a�]$t(Sk��%�f�=oN�f�$��#B�KJ�Ȓ�����RK�N��^�?��z��<����<ߵ��m����iH�Be��y k^?)���f�sKW_Pv�@�g��l�&%��㋖C="p��^�<���W���.	Ix{����n~Q����12�v���c�lH@¶wy(1��K`�<$�N\���Yr+x�