XlxV64EB    1800     850^���Z��6�_�7�� E�'d�A
V��_oDɋ7u�k�^� ;��O�wԾ
A�<������l���\H�#���l�|�Z��.Z��rk���1�,�2ERF{4���Fݢ/,lզ^��V�]YD�g�ҋ+��n�t�M��m�;�z9����Ւ�;��{(Ew�+��7�Ɣ�&�	Ʌ)�6�A�S*�'�褧�[�-����aXM�z0$�4��`�̯��� {�F�WIί(���8��b#3F� �3ρi&Ƨ[��5�F>4�W��m��λ���N߆�v�x�e|N�vG��E}(���pF2�_�ȋ���ĮKN�%�7�t�@�ډ��iT	��G����׿�3wH7/��W�Y�!A�t3�H����H����������TD8WF~Z�#f�����L�[����U�ޭ�;���ˁu���K�~`%�,8��<u��G�6��C4���;��!��e�9�:a^?�?hB�=��Q����-�sȜ��������^���
���t�us���Ic����tR��$�O}:3�Lǂ<�V��|)Oe;V��r�0_u߃I͉���g�R���]&E~}srGo�jK�����1�yԂ��Hg��^3��k�]wI1�	�5gF
���u�ǃ���/`��K�0bв%�%}q��_č�����أFK��-~»�/���0����[�C2�)�J�1�9A�ԩx>|�nY�����mj<�����_�8{�8%/�=�vM���9����B�Mm���hpΔ��nW$N���f�h!�T�G�wW�K���t�Z��o௸��A}��_D猍u{�����I�#�xUڊ����j�q��3�gj�S�U�,I����&�haO�����~�|�8��1�EF������(u��N����8>G��M�MϾ��� �';�V����	��L5[�?�$�(A�{Aw��0�⣳����y�k�ܨD�[�s�i����٤�u��Z��]�g�%_����iSF�Πz��1Φ���F!�����<���Hp��f¤������A&���ȡpmY���Y{��[��׹�R�r���u�ć>��.�TO�#:��X���P!<�lR�&�&d+|I^vU�C-�����@��F냃UV��g�Y�i��"a��ʆ=�>����)� "bS/'L?��.#	�׃lS#_ f����r-�q�6
�=NMT��橬�j��c�����^ٚ00���ϸ�-��.�G@�o��۳�@���ܲ�p��	lI^�*�	$�V����Д�i��e���^�I#S�ǪS	OR�FSU�o����x�U4|�|��B�f�	����L���P���͋B�?Y�9�|B�?@�Q(�foVz��6^�� ���,�uj�"}[��;��a���"�8�)gl�f����+��TX���6�D�"�������]i�����~09-��]�b����B������-�F	5��h[��mz�!`fy�9=LleRL��z�󡕚��u X{���c,hBs'�2
�x	�%����ɋ�O<��T3K�^��R���'**An�{���I���${�����d�w�sx��c���ٿ ��e_r9��XT��÷ɦ$���ut�+�.�A��m���I�=��j���dg�=��X�bϤp�]'�,;������pT-�X�o���Z#V!n��q<������H��̤��zud\|3����T��\jd��G�U��G�8Y��T�C�� K���{�HD��k ��,��'8x��mj�'����|}�(���nl ���H�W�f�\�^/�BˎV�3ل�����"ʁw�޴��ڃl���z�H��]� �p�Qݢ_7���~���0�K�3d��{�x�L��Y��Ph���@Tn��:L~S�e����5K;^)\��g��\�%I#mQbQ�����k��:�y�A��S�dF�t<���	(3E�yR��i�>�����+�(���p2��)�=�]�"-�HZ�n\��D���;��~Lȶ	��viȶ	V
�a�C8@vq�D��.�i�2�����L&��b�	>�