XlxV64EB    8378    1e40�Q��ڐ�,�R�B!��Yn�d�J�1�)��� FR�:M�����J�
�l��l�6�@OW���E_��h����cF��R�ZƑ�cST>B��@u�����-b���g�ֻ��1�w7��b��rX_�������P�R����.c�N�7���^*]J�!�� �g(�Ӑъk��(��c��' �)���%H(��,�5B�4j�Na�?Ӥ�һ��P��80	�yW���@#�&�Ջ��聲��m��K���D�b�S�=%E!������>h�����܅:;ҠVt.��1Þ���J,�g���
�E�f%���u�� �CIEz��b~�t��!��7t��H���o�G���~P�iek��͸�e���w>���k���f�]�L�j��4�;�Owi7����v�w;�ҁ�:#�Y��w��,���
�:�}���(���s@,{�X�����C��<t��m���#���khq	��F`�VT
G!v��b[���e5ٍW>�j�q&�:�/�b9�R���?��-�'3�r��	�ؼe�F�J����?��-����I��Ճ/�4�k�G3b��p�=Z�{D&�_�����47Ż�o��?�9�H�j%kǟjG��s'��U橚�N���F8�5�_�	tq,�\�
��,A�o��)_9)�\g�L^1���S����E�е��p�>���j�X�BR�h�� ���7��_��|?1 ��,�P:�4H0L�������/o��KdL�f�i�+-�%2���uh��D{���&A\�~��k�~��$i��� ��rH-X.I�M�W&����H�_9�P��_��s���N�U;K)��ĘX\�iY@	�L��D�Xzz�KR��NK�&;$�D&9;��7�Ë�߲���*Ѱ�.�7Tb�K��l��`1��W������I�j§8.k�a���Q��>�X�v��e���5�����RfA���(=���T&��KG�|�Ҕ'�OUrm�r##O���5T��7h���������F�f�dn��.~�C�3��*���9FE�7渞&��i"��4s�)>��v�M9��D�Yc����֦�':��^nf��D�DQXY��G�F[5o܂t�xJLݞN����Z��t�um��E��}u,����2@m����K��`���-�,���|�Dy�t�bb��/	#���͝+w#q2��6h����{)�����Ȍ���nQ1*a�r����"�*���Q�t%���aT2�W��+C���z4���iL��,�`�5�Hkk�A��eM������jD�q��T�R���=�U?�{�zZ�H�0�K�Ƿ����|���1���Q0:z���责+��{���F���TxyI7��a���SW+p�m�M��d��k�gk���6��M_l3�k��q��J4� ��r�(�t֖��.Xی�k�u�u��,�X�	�%�X�,-=�n5�&$��>���q�Y�91͚D�1ٖ�!��Z�R+�&M���U�-� -�����Z���l���L�RD��>���3���M�&b\K���K��!��'}��ht�����6;��<c�Ә��Y56Or��zt���տ���i��?�7�+J�5���-���Y�ӿ�������s�����"��_IA7�����@;�
_@��Nǁ�o�C��@�hH�~-���&��0�{��QJ��h�\;>k$]J�Rq���)��k\.�b!���̧��&B��3��~��$J\$5i�zWC�M&GB������0���K�	�3��.+�+��J�t�m�������&X�ߋ-q<p���zm���Y���A��rB��ך�� H��>-�55!��P�S[�*N�F�/��B��;�?,��PG#�_�g8;Ve_J&���~�hY�Ĕ�1U���u�2{ƯWIrA���Ѐ����A8�#d�e���͌�;�	�<Ƈ����D�F�9�p��9F��o
[,���أ�>i��Q)����b�# U���f񺡩������,8��1k��g�ENҨr}�i��>v!wJ��>+� r�L���2�g_����n��W�Uh~
��plY����Q�iϮX
�X������@��uG|�&c�P�M:E�`�(L2�0p�hr`B8pXK��&yp���/<���p���)����˞ ��C~�9����P�ۡi��z~ٺ�Mz��?�8n�C#���׀4<*�	k��p����Jӥ��==�l֥��C����v�w,��^�YM�K��|�vq��A��� y�bw���E"H
��B?1gm�C���ӎ��X��ݣ떛�ILZVE,��ͱ�N�J��9���	�)ֹY`����q2I�S!N�ph�� ��.���qhD�,Lz�A!�$����/:q6y�	�e5lc�es!���O��QD�{�d/�c�b���Ґ3�oovP�0�Hp���^��Z(~�XMO�v�Vi��0�2��e?�T  �,YF�5_  �_֦{�=v"F �z�qBL�:9?��T+'�u�jṆ�Y]��f��}MK��\�,�l^��1��(^!4m9�?�����'�~����^#�
p����il$���[À"����ɟ�U�0s��F���2��n�;e7��1OO},#o��'�r���?��%�*���i$#Dޘ��cM�S�@��裍�I�?��Ⱦd�����MP{$o�$�h"�?q������ 1+�Hr~(u�q�DDDW���H�b��f���ڂ���؛©観hy�8s�k�w��l�W�;���d
���B����YU891��D950�S�� �8��(�顁��C/8�۠ܪ�j۽��Ռ7t��� ��5�D.K���=z�H�F�q�JS?��t���N˖lh�S�Л	�"{eν�P�����w�_�����ߺ=� 5�"S��;ÅH"��U���&���Q��6 ��y-�ը��&�FG�8�^d����@ܬo]x�I��ï�_�٧_�3by5|�Y��e�f���U$�p3&'8�ԝ�'��������!������B�1t�Ӡ���֝w�	j?K�u��.~q=<�G�,*��YO�-?��,��ZW=͆D�6V޼�}N�3r�p��Yr�]�n���\��G��㵩�� &xD����eUN��ā���)־MÝҜ�
@�͏H)�_�=YPJt�JLkш�����i�D*��dr��H��YĢ�$0."2��$:~��2_6�o�����($�){Mxm��$i\�a�`҆�� ��"⎔6�ч��0u0\E�<�T�M�����������Ax��/>��g�q��9�B b2_���h�����jS�]�J����69�ˮ��M�x?�����CV��������P9V��{/�o�i���ڲ�f�8���/Hd�N�ŏX)��=H�2�g��LB�_��#�%k�Ng=�U��ݘ��.6dʹ��|�<�5"<d�w�mg��f�s�I��2;۩�s)D)6����[H�T����l}b���=�H0��[s��7���{t��?#�iO�!z&~���ʣ�yN�p{�o��}1�l^�@TB�N�i��_�x�� ���5>V��?���e�<V��v��L�&�be�ȉ��z��A��&��^�8k�mR�t�ua����Ef��7v�9ES ����n�^UD`����AX�f�L�zp%���%@P
Ɏ\ى��e���MU��)�@��6���9�T�����/O��NA�#��^'�$be[Y�nZԆ2f>z ������&�`6�XMA��Yv%�;N�S�A/+ha(�$��Pj��Q�@���j�(r>�� ��Pn�:w�y e&NCE�W���K���= 1�+�����?2{��Ϋ�G�MI_���|�ԏ4��_�(<���J@�������2�i���>K�D�^��g�Jx!���u<�#%�?ӸlyJ\�'����D��R����GN�qym�Ns���'�h
���@4���H�lE`�$H�)'m���ž�e3v�b��f�)�,V��������c ��R���ȴ�-g�s�qʹ=
�\0���SȎRa�)|��ɂ�FL��
���\�bg�j�-d+�#���,�����J�G�ç]�Y���k?��'룄�����"��E�.��������j����&�2|S�M��������j���.��@L�{w��3�w�l�9C�6\ݹ��u������@�UŨwv�3Ӭ�:�S�Eq� k��r�_f�����P�W��l��L_�C�
0���L���9�IaDR.5� .5s�8��X�Qfn�~���Wik��O�U�Fa���h�$��b���VQ���-@͈��{]	�@�aƩ �\w��qka�r)6>�nL`�)o��w�.�ᇹX"����#Z�M쫃��ønS	�>A�9�ʆ�g�h�ӂV��n7��H���8�\��������-��+��͡�����ѝ�V"k!�ks&-���2[^�u�#{��aa|eφ��o��®R����� �m.��G���|J��N�x� ���.twl��E>�������Rb�UZ٥W;�\Q+̅f�{'�|�V�Vsi������"E�	��jV��-�Aqx%���, �TR\�E$W�X�Z��ɯ��RG��vKN0C'@y�DI�\^��'N��D��Ϊ|0�,>�C�{�\!��a�T�WK�(ߝз\�LcR�j��w�٠k��P4ǻ+�$Y	0Zu���2ό��ThV���ͦM
� }�.a;�_f.�\�L�V��
M����o%��^n~!`:γ{lG�]������}mY��â�ak��DI�?}h�:�4�j�*��1+�[dLm,�u��b��V]�� �!DCc3�Q�,�J�bW�<Ͱ��4�Q/-aI9e��(]�v"� ���!���%.�bvYKT�J��q7"�A�C\�vJ�&�j�C�b;���x�ѯ����׮�-��ɾ%}ǽ�.܆%�ʣo�1U����(E��ئ�i���D/�I���)v�$πr��L������y�ބ����σ������8�Ux�Xg��P���5�Pb~���Qq��N.�����K��G8=g��z�w��5��>mHx$�r���� �[�Tʃ�=oK�
���1x��h��E)�Z���7���6�'�oI��
ꮮD�5ز���%���<�w�-1�0���W�T��\Ӑ�L�P�3�;WT��������2Z�]G7=}*�b������443���yWq�5m��ǿ���~��-述M�	�=s��U�_�����h�t���GU��s"*��;��$��1�WI�oï�>2�c7?�>��O&��?�d�T�+?��D�f��8Y�;�@�0�.K�@��r������`%��<ͥ4	6&`����~�n�8��!�P笝�C�p�w���d����������� ���G��K,� 9U��F��͢�fX�\&����~���HI��X�l�	�R
�[Q�S��R�"��U6�0,�G�YL$X�*��"�'<��ǟͫkT��y9�a�U�Ľ�ߺ�"aF���o�c�.��MLCyBX��=����vc�^g�o7dq16�ѐ��6?��@��PO{/���I�i�1 H���7����7"o:�CػV3p�I̜J-L¾���3��j���������3�<\�+H�&�'~j��d,
����k����3��%���Ͼ[l�M���+R��U�渀�A3S��x��ۗ����U�pG���<_1r���������L��qb疠q�hb��b�I��/K��1Fl�����|���-�������g�@l朏s�ϭ9��Q�U�/������J1ΒEZ(2�����(8��2�O��$(C��� �t휩G�E�9y� .٧P��u�}�K"�C�A��څ?=e����k/��p�OR�<�A&pf<�1�U���Ò�"�*Kթ� ��2����U�c@��(궯Q������j�Gz����tQ�/_	8��Y	��fѱ��z�BZWވ��0�k��/x� �&v��L/��N����*���4���X�Ki~fk�1�^T�Eѽ:�2�2��J����s�J��ENE=�:�!�4��v:��1?����F:��4*L�ɛ���X=�&��)޺�PJ���� qG�5/��维����/�Ю����D¼:�+���{Q�HB2���A�]tc���˓��Y0\{*��5��̺�(ް�Q�yƬpRH(A�n�����%�������O��0�0|��LY.`B��Tj�f�B��XP��Lz���8�	��)W��ա��v݁
n�X,H?���7���!�'����5D}�=���F�@O�j�R;ʲ�'{��w!c��X Q�
�P&�D�.�A����,�F�<EQ�3*M|�����#�����P�"J}�lH�%�-�@�ky�W7������hç��C�� �^��2/
Kӄ�`jEeي&Ľ�F�&����N/��%�1Fi�	~�ڌ��-��.��ik2��Z0-�)�C�_�[y�cO2��;Vi-��k�vL�������N��?��[�ɥ�Q�~<��e ��XI~�ŝ�9�n7y��#6��(�������ރ�Ԝ&h�&�
�����v�I�q���חaˠ���c�I�1�)�F����1����p9�<�[;)\En,����� ��kt�:h\�kZ��T�Cn��|Q��j��[����l�e�9�CP��Ր�K!gm�u&"؝ֶ��'�%2�Tҕ�P�V� �֞4���K);�E����Q!Ge�!^���Di����ቍ�8V얹L���	�]�􍆥J�>V{��9�ޯ|���;��⚅�j�ə�bj�+��$�D��U�Bg�I3�a����vqv،�hQz%c�k��<��+�a� ��2X��ޙMg�&�ԬΒ�B��?��`;zV�1q����F�߄��S](H���h6lg_���0A�-N -�'"�y˒�E�N5�D���Ǜ�v�0W~D�b՝�2�a��/]�u��Yu��L�K�'�>���g�rD%"\�6S�ݞ���Y(L'׏P���W��|K�N`��Sk�!��溶BU$�}ُ��wE�s��F��jz1վ�B�,&p�@�s�eB�Z|�P�����%��bI�C*�V~^�bxs�pz;��s��z��@������fA�,�Pޱ^���(o����p��rtϢ5����s��̉�����2ϡ �Q����u��a�e$Dӡ�E�Q��J�[�_�W8�-�1��h3��e/��x�Ʃoԡl[���ݸZ�z$#�L�;D>�������`���Z�=^�]|Ə�|fX|�z���0R<�v��6i,0)�O6�=�G3P�܇��~��5��u���S�DQ7�0f�+#������|J��M�-IBB��7��4�$g�i�F�n��Lg�e��V��8}�٣��������e"���Bփ5�YZ�)�e�cO)�A=c�wp��-���7!�G�Kp�R�j�