XlxV64EB    201e     980Y��D�AU�ѯ|�-m����,��t^&�q���,�{��m�Z������q~S$�ڨ'Ae���~�#�� R�iU��/��R`{h#"=���3��D7��X͋�6�8�S}͂W����f�N:��iU�(�]j>�Ar�H��6��Q^���Fp�E*Μ�_�W��N��6���3q��C/��(^e��U�Q-Wf��f�PG1����'������YZ���������:���(��ۻ1˻ri �6V�=���� ����6鈜�����ͣ��v��2�}�9U��p�8`� �v�m���Y��M�Q�+�w�T�U�qfOdEJ���8Q|�3�>�F{BcB?v���tM���&�t�Xu�{O�k��~0�.�}����3h\(Vk���W�{ ������ܺ�������� ���f�Dx�j�]�F3�sCD)Au�t�'$�N"���)_znw�ݔ-�۠.D򦑛�&��՞�1)EV��I�zb�m��/l��j�j']o��X�c4��\B_�'zI��$0	zsA�
2
����KJs�_F{`Xۇ���8���Yo���t��&o%�3�-�7R��"WUzh�/`H�>�8~t��Yo��Gv�.Z��j���20o/��ܤ���f3�.�!���ܺo�D߃�TI�Wz_#.
LM	˄�`�QAbl�6�8˗rP��}�Owj��kӋ?�~��2�ϟ�s9�3�yq��D� 1�zo٢�;5�g�
��L-Hk�w�����q��WR �b����R���q���=��MS� ��Q���8���� �օ�i,�,�M������s�L��?t��������^'L����aߛ�c�C/E~�<TRv��8�!��T�	���P�N�QY�I':ӽ��h�a�����Y��(���̄�.��n/��O*�9;�:�p�;p����9����Xk� )���w�Q��-={\�9d����}ڗ�U�����SL|�n��Y�B��>�NW&�( �s#'���&@����B�V��M�kݔ�_/�	��o���hABqG�k�dP����G�]t�	����ۜ�>P��G���ĄU�h�:1Ճg%���[7ʘhu�C�al@啉�������j��]�ѧQ����1(��@[��4-���X\�Ę?ōl.ؠ�P��
^w����^c��W`�+�<��^!j;��Y��k��[7�e|� v_Pǌ��H�}E�E������'��!�)a�l��ؕhղB�/�L�0�z����ȭ��Ļ�������e2d�o3�rZP7��7n(���m%��b��o��X#?`O��;�ͧ/D��@�w����Ӹh�b��>�8��K����/4��7=9�" �rz��gTӼ�葞O�Rn�1���~�����C��Ã�u�'���]�<�e�����c�"nF�$��
�y�88�ѷd�̗��$!#^�����~4��˼����$�˃��� 6P�'���Q5/�ݼ �B���"�� ��c�"O��[�UPV�x���0-1�k:f�%^Y�@o��ʤ-L�N4{V���;�X/}n���ZA5���uBӻ�,O;��Z͸��vp���ޭ׿��(E���
 ���`f�C�Oo|~QѬc��1N��[����[Q�G�7hڟxgV~���\���7��a)�8�:�޾	׸*=T��f�KF��0 �m�}Z�*8��齾�k�ly^�㞋 ��D��Y����� E���Ջ���q�P�"��%�/v�OJ�����i�`�b3���0隆y�J̲���;��h��`Qɴ����A��ح6�WtOI��GݤPΕ��'Ĵ-��>�}Ȱ�L��Z~��GȤ�|F�Ru	��u`Cx����1:�s����[ч�Fʂ��@�)Sk6M�(8rc�pSus����?x*JY{�-�`��{�� �By��O��K�]�Ox��klU���������%=!v"�I��>ɤ�CN���&H%c�(�{��6����G�� i'� �~+�c�Q��4] D"�x�d/��%���4�}4��U�!59Mm	�0���y�v�U���eTmJ��UV06��*��Ig�(?g
jW�9'�]�R�P�-��-�9��A�(�?+k$�+:E�(�/���?���-OD��v�_�~�%����G�m��ъ�8��/�^���
(�������½F�|V���{:�*���U��PEw�i+��R�ů3� 0�}u	X#sn����{��p7pհz�*�����OrH�Z��HfVIA�}4"��ض14fYz�v37iG�Tg��}4]:z���U�W{g#}�+^�-��5��0r}lre3��~�2�����/�Q�`�iCg2��)Z�K�[x�