XlxV64EB    52f0    1190@1�5��k>�I�؆�yB'ne��
�o��A��\�S�]�K�d5w�Я+;c'X�i�o��1Ѱy���{!�}��I��,����gA�
2�Μٮ&Wa����ܤ+3��0�V�?M��n��6]!S7�1?ӑD3bX�ɮ��8'����f�Oѵ'��+;4z���| iZU�垘��d$�\�(��=��sp:��#A���w �Ό�G�E	����C����hK������`�o��<�Jgɭ�X<�Q�e��W`�T,� �q�[4�^��~��.���U��tߑdIiJr�s�Yn$��`D�I?y��B��)�z[t{6Ժi�ʈh狮p#
�� �?������ȑEj^d�ͪ$�A��aBWW��g��C=�RRA����ĳa�42v�W%���X��҉�J�, �P��)Lsp�Y�}��ʶ�����Ӆ6KR<�}�8|>�Vm��7n����=K�7�~?ʱ��ߤRs����(�8���z hI�&�;�q}�s�f��a��΂���W� Ms�t#�Mf����U7�E�O�kg�V�B,�G��3��Z'�����x���讦%P�
��[n��K����η{�8��*j,l���~d_E|���l-ɝͬ�.�i��ũ��'v �OE(�V�����p��_չO#��AoٯK^N^:�u�S�ϑ4)�#4n��8qM=�Z��|���'���r�����ι��P��8P��k���`�m��v���Oq�O�uo���N]�{�/;^�C�9��6�)^�(�9Xo���|���f�z� R	
;4^JR��+��t-]�~�	���e�!g��v��AiYc�r %L�x ٬�[�'[b{t�q߼2b��2���y��6�˵NŇM]�ƶnl�o��(c���N%�R�T��XC�w�̢}�c���d�F����M�'��Y�v���a(�w����{�+Yw]i�i��	&�$
k�9�p��2����R��C]�2�,h�$>|8�����ԩ3�Y�4�ZDl���T�D�@{T��8
�!�H%B+�2��+�xf�?��U��$_�"��E�S5��_K�c�Ů[���3�(q���X��I�ƅJ
��hh%���#�h�`�+<�z�벣�I�,bniK��g���̼�3�웙�-"�ۥ>k�}��):)�<�)�8`���ӝ@[���KU�Z�j����t��Sy��H m��䄷9����9�=օ�v�C+^��Mac�ѿ����O~�l����ƙ@9p�͓��YAvc/�r�N�oW;(�lvL�Yw@QP9��ȋgC�CF4���#<#b�kVl>�(��ɒuL���G���L��k&�ϭ�L��Y����%ٕP��ivmZ_�r��j�-V�����W�bӎp!����o��$W,*��
XB��\J�T��\@P��?�E���J��N��r?E�������>�5�|�G��ʺ/���gU�U�3�sSD>�-����=������r�s��ps��[G�W�ۗ���FÕH��b[�մ=ԙ���1]��
���#��I��7 �	�ۛϷ�8�~�[2��ڴIx��-@"��G��.�T��:��7��Q��j�����k'/����w�g���O\Z=8L�ad�[nt~�0SB�	�:�+,Q�j�-t�
������}�$TDqE[�I���;��wV �r��cNj�܂g[ː�7i4E��O�g��Nm�j1��S	ݵ�=4��4̖�5$�V;[�4��t��JC�e��!��(s����?J�6���Q�����~۬��R�y��I�Q�5}�}�ee�N���?QE�������ۨ�H��z���Pg�}ԡ�;�&�Op� {�l?Of{CE��D�I�^I�@�H�(�H�w�s�`��ƹ��s��I��{Xsl�rU.�Q���E�����ߢB�B<`!*�5r3��L9lԐ ��7���&2k'y�T�����5�Ϣ�����S����H�H���eRt�֛룆�ĕK������u�@�*7cO?@�F�0���H�/k����L��yc�#�O_L�d\CP�I?@|��X3)`a�\��Nj�`D�==SR���#w��2�Bh#A��p	�~��oR�p��)#t9����G���0�*��k�J��p��N�{Mɫ�y���_�7B�Xvq�6�"[�u�\����W{���n͑[��p��HE����9=I��ɇyn���|�^I�C�7�e�.]j�*�d~޷\g7��F$�j��g�a�����a3�!8�,t|�L��*���ߒ��Ŵ�KՃF���=5 +�\:A�"�@�8�z�Ǩ�N���e���֦p.�9Iێ�í[���a(@���d�"\U��@����'���t�fGG3�vNG@�)�d\����v���� ��t��ͺ	��31�⊈��7�P��@!B3
 hxoL���i��RT�&�>c��̢�=S���M�#R�~7�}����6����3i\J��G��u9i�'#�YRj�ۨ]E��4�}2%����a%|G�0{�A�6�����!"�/��I���i OA{%������A,��1�U�h�RJz~����n��<iGo�z�f:@p�\�)�_�	
�8��O&��҉�&(�(+b�_�@S���,�K��!�S`sr�2���Y�q>���E鍭�_���:��}�\�ڥ?��{F5N3	�Ve�Zͽ{�yN9�9���	���Y�6�W[����3�g�p�\`�]U�E��S����<����'J���w%��kn�ax�W=sF�|���\�>��37q�Ɇ���u���&p�`Qm��a�����GR'�,�#�q�}�1��j<W$���/.lja]���Q�����
`mj�(�����h����N��O�rxmq^x.z���5�6��YU��ꯂ�4�
�_sh�����$;]�M����q�K��<�4*]�j�q)	�����%���s�le[5��U3݊��Y��1�0y%8�¶���O�ȅ����U�rC1�D]Bp������fO��;�_w�gÒ)��k?����L6R��lZ�ء|�ㇿ��w4U�	"���k�װ*�������g�K%��8J�
) �}����!7b��0�]�KS��Ĥ�t4�7���s�!��?�K�l�@9�VDx?h:���c0�ioﭏ�8�uq�jy�	�l��T�e0\�)�ǎ�E$z~G�=G̸�ַJg+��A�^) ��.5�D3o����a�o�A��� GJ���ȫzh<���l��i�!��Y�y��pC�Y�'�����PS/��X�%�+P�=�Dc�r�d��>q<K!o���L<0Ք��NµZǷ��:	~�NP��Y������개�*�ɿ��һ��0�q9$	�/��,����H���l�2��N��?�>�HKX��N 絩�[�W�b��y���:�/nXA'�Y�.K�1��!���j�ΰ����J�:�E�T��P]J[v��%�����H��2����cߑ�R8��gV�������bE�?z.%&���Z�?�'�c�^�*g�+Rz��

]$��`�\�t�E@uc�*�P>[[,8YoV�I��&$�h��}��*�D�-����X��'�SQ�X���^�B���D"3�ŗb(��|=�	=�8�����>d� �������:]��-$vu��>�94�=���$����;V��Z'�D����;�5�f�ve�UeL�
v���mW�tc.�:@h7�E@���۬���Yϸ/V�ꈽ�]�0�^�������Ǒ*˔B@(�mɉvua�:R+��b�)y�T�����HC��k����̑f]0E&��q��حXw� ��j��,筲ј�����L-�ݚ����ֳ5ذ
�=����+s22Lh�>L���N�D'-,{/��P_V�gj��T���8R�x�ݮ��r���|@"��G6����dY�-�Q��ux^0�=���ނ���Ssj�����υ���+�(���T��ܑ'n��)\,���C�  o�Wk8Nw��9���Xס����@���U4�2��Ns�۩.ֆ�)�뺴��l�tȮ�ҵ����֑�8�UfCchy|�gv��?N�;�ٟi���9��ɑH'�*C�S�2��)�N���M�+��j`�<�V6C��᧞&���M�X���T,���w�^�[C�\WF7������]7�P=��!����
�b��R�(��f��(�{A�5cM2sX��ǔ�g��ɾ����F����h:��&���tp/����~��N�A�.��D0�x�w?�L(#����W�^��y*�<h����KSvIV�Щ�B�	����+<�<�%����9F4\�UDD�ڄ��^+`��]�CJ���mw�K|,�D�m���W