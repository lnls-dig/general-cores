XlxV64EB    1d57     9e0����P���$�.
045<�l ��|'c&��-@W&�C ����Y6.��7W��%���Y�-�.�� �ف6�>7��ӿ�?r�&�r�Y�ِD��JmF۴�AE�o��ϐ�%�ȅR�+�5(�i9Au���v�]��Ƀ���Fy&�����"t;�h��r�:���b*"����ʯ/��ٲ��X��� rS�����&���6�0o�Q^��f�]E��N��,+�~�\�LR]d�}R�H��<^�F������F�9MN��T�*MBX�8�L������y��9�kJ*��M45&]�'�o޿l��@i�H�Qل�Ϳ|.�9�tP^1 �F�k}�ׅ�YK^����>�B��~��RhJ�Z��~)@^!�׉y��P�g�q�vD� �$�䍨`��"Y�W�3�,�2J�}�$A~�~�S���{��� �Kէ�m�A,�x�S��[ ��$�Pm���� �w?YY��E�E2�Uwa�I(90� !s��jD�by\�BZV��]j=�q�_��.��N����y�����a���ާ�������a'hEE$��"j���iMiVYWCJe�9(W&�|����-��M��LT�0RTϊ�+#�/�i�jA3�9������'�4ۇ���d���ZkO�QDI�#�\z�ώIg�>r��r��Q:�o1LֵNl��:�W������֔�Ս�`2c��!����=��})�b-��b'Z��}�G����I&AF�:'8��,CsPj�<���>�V4�C���]L�VM��NT6[���K/K%�?�!���ǮH��l�-`}�W�Xo����Q/z�k��x,����|�O���]���j�U(�"��ğ�:Ҷb��',�֑[so�[�'�@C9\&��_Lu�ږb�@d�P�1��f�35c��LO�S�\�IN�;lGq'���f\w���QU�V�&��~��`�$,p�q�L\FY�����\�6�(�� �.;Ÿg��}�N����@/9�\ZL\a-�p�@����v� i�53�`X�D�:g=�w�`�c��e"s��Ub趃nCNw����]�-́�8�.Zږ|�)�/,	F]��W��ށ�R<�wc��{�������yJ�!t�-5�J�����ާ��m�;6��:B�3pC��&95�)�M6@����O�bK_a�- ����Eu#����[t�||DpEۈ;����`�#�[jP��%�d�(���\��r���U�9Z�JV+ *:S�/*ꂍ�V�ο�C����.�ռ8q�w�c\�[�R~�@�/E��?����~I^�Z���~�d��h���c��:�B�/�L�x�PmO�C���Ez)&�)����H��jcY�n�Z?����>B}���y�.��2���#��Y� `�'I�'k�E8&aUK��UV�t��QR��*�o �-�TS~M�Qa$ԑx
�M�����(���ϕ�_�˙����	�"���t?�4���߷��x0U�K���)5�l�Ǻ�P?)ަ;3��y��
3� ���)�j�n�5�!��5V�6��'yR�D暊��'���^n�'|���n�2X0��	��@����l�"`t�$���т���$�#g�����F���嗮w��QmI?[0S}�&&�Z:��&�
-hB
k�Ѝ�-)ԙaTl���
 T�А:v�;�Ey�G&2x��]��om���A\��8�����uo����-��F�b������jJFE���p1�SlgP�,L��C�~��ر	��~dܥmV<��-�5� e�}w���2�y�J`��]�*�ɀ���om����?�K��7�\�ɣ�����9/�R�Ö��V%��b�[4��ͨ���y��Dh��%u����)F>���
�u:O��'>8�!6~�YT�	�Eǚy0ҶǫR"7�&������Py�ՠ+?Jם��j�Ï//N����� ��V�h�)�*�7r,-���aS���~):#���ԫ~8��ɵ̝fE�t�v{ �{X�KB��G����gE�&�x��Em�?l���H#��t�ַS��$�a�1h�JT��?x��g�pH!��KL�	���1M���]�M��<8�^��	|������@�N���4��y����a:.�xk֌��@3�:��Kb�"���}o���A�u�0H􄻠�Y�ح��拉�+��`.Pm���v�u̟���"R)�FS�h�ѳ�*�d���?J:5��5Q���g�S�[�C��yy��T����OUP�b�_/vҙ�g87������Q�#�����Z����ZUͥ���.��s�� �Z1��mvyY����I����7[����ˬ�H���jm�F�*��y�6���� �c�H$z�FJԞA����ݤBCY�G��so�Yj���4��[�c�k����:�οjሮa!r��fΪ=*QG���: �]���{�'R��Bţ�q��5E�m���S��