XlxV64EB    2707     a80��d٠�8�
�f8J6R4����u<*�^������X_�>���O����/I�a0{D�j�x˘����o����b�ͽ!�˚�P�\�_%>���o�$Nq���Ek�;�X��/4ߓ�h�@20��zv|�A��dE|�'�!��d���!�e�F4���ܸ����u�BN`1��a�KGf��>X�}z2An֬��fRI�Y/<�k��I�M��Y�&Hd]��N�z���o����S�s�"�]8��C�6�ǱZI����vgH�ĸH�c����($7��� �c�ѻ�����z�D-v,^�0	�T�q\��5ڶ1��)�4�R�~�7���ɳ�{�ڛ�P�Ö�m2��o�s��jA��	��8�?�	1����9�0V�k.+��5�~}A�Ԁf��$��o��D�J~�u�IoO�0?���_օ�Gk~��9ƆD�S���
t�� �����Fov�v6��L�.
P �Rq�t�����h��~�]lvؠ��x.��i{�k��Ѽ�I�	�����:贫&�?A�G�:r�� s���:�c��̀`:Ȳ�IR�16��*�vA��	�JSQD���:>闵@cSx�Vg�v�P+05�!hl��yÉt:c��R����`V�A�R*��;h��~��: ����;���J���N@H���D�<ٸ����FM0ح&?�Ap��3Q��WB�|U��U�1Q���Z^�a��ώ~WV>%	�Y ,񼏵ӱ��9ڊK�뀇+\��R�W��Y�7�O�ƍ�>���q�����,k���vU�&��g�	�/�ZNg<4�L��L�(����}�}]�<hl���d`~7���Ę�Bgg�����Ft����	'��G���<z�H�[��M�_���@���jU�O�;�)Q{잉�-b����^cgsRE�!,�2����oxd�jj��~����u�=�A%�1�uN�5H� \�?lMh\��z�'|p�}���ŷo\�=F`I:%��:���$�:o���U��*�±}�b�!&ŗ����^j�>�K�%Z��*�����Vt�9��{E�Ӧ�F�	�,���ʿ���n�8I�.o�S�Pk�r����ik�'#��+�"Q�!kxe�j>��$s�^)���L/���]�����WҀ	�dX�D�_�����T��TC+aʃ֏#D���kcX�ćP�!�G�6�bʪ�θ�ۮ�������(�11/g�Y�}�H\�K�X��ˍF\=?��{V#J���\�r�d*�_F��'5H5��.��R�����i���f��;V\��p˧�j�1���V25�z=���@s�� ���;a�
]58�9�V|ى�����Mi�*+�YZ���+���ۢ�r�6�
�8���et0%��巼>����Լ�(��Qx�Z`�~�1�Q��q���O">UU�L������nk|��gm.o�lawJ�!*��מ'�nEҟU���݄�	6]��v3��\����4����=]�3R�ڌ�aL�'Oı��-~F� 3���Ǚ�W ��Ae@.)�굢XA���o�J��C%�V��H���b4)JB��@!]n~�=͐F0���zs�d��%)F>׈��a+�q������J��H�N'
uÉ?�Xcْ��f�i��P��t��7l�)�"�>m��/�M� >4�xQU�\6�r	��g;�<6O�3�ҡ���ǂ��2�,\���Ze�/�U"�uE�����P6�k�{���םf�BH�7��f�!��#�L��� �N���.��=|3��̣��'�*�Ĕjq�^��@9�?�@����@J��v���LrS���%ﻲx�cLB9CNtg��ʧ��䵫���؇�UQ[�Q$���-��#oX�pcOT�h��I����.\
`�8қ)��=�
Er$��1�v;9�U�w8+��#b�z��Q>�%�	�JJN�6�f�׿	�׻Ί��/�I4�4�3�`_�O�э.��ޅ:oͪ�fZ�+2��HiH���n,�^ܡx��В��40�m�o��tD/� ��'�!��ҬV�MXs���Y�*%00��1��?A�v�|�����0��W����k�����n_��g���� ��x�΢��[E�A�Ő�/֫��ʒ�^��j)���yw�P��B"�W�F���+�7�O�ys�����й����|d�!h���@�������`���|��Xp�,P�fs&V=��7���_)�"�\7�Ř5���I�G%	[�&�w���W׿?0&��� �Gg؇[J&��&�׊㩟�7��
i�O��X�C[�9�Dqz�]M�ǽ����G�2�h߱��U7<�� ޅ�cm�����]I}��r�@q�*�Q]U� ���W���xHV8f�e<i��-�19J'%{DR/�+��aH�0)M�
dSe_.ؒOf)P�:���}YB�z��ڄ�
� #ȕ����t��$sً�
mh�I9H�v�ԧ�	|G�Yd8B���H�;�a��#�����H<��ȋ���qj���}��OH�W�������W=�2�h�AV;; �_H"9��"�K����㆘�t�oҶ����I:!S$��N
�>�4_&??�Ȕ���l󿔗�����q}�)�ZX"