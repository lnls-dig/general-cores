XlxV64EB    5829     ed0����y�Pp��_{�0و9�^���[�o�٢��!��>��5�h�j�zl$�y=�A�X��M��jF/���;��+t�@�KG}P�����ێ'_��h����&L�÷**�1A�:���9�q,�� N�զRs�F�i����яdHB7#"��a)����`����@�1ƽ�e��8 �%�vw�����I"�s�Z���E��1�(�p	�y�������e���I�X���8�<��!����7s���\{~��J#>S@4%r���������Sz����<��/W��SǑ���jv :Yb�!*�/M��a4�b�����QnH��7S^�N�V��_���&N���v�lg�K����ҁK�@T�w����w�4��Y���	�&M1�LF�JZ�9]1 �L����Z~�*CH�x~�Y����$��X��F<5:;��,4E����=ie��8��H0/g��=T8:`�"<��a�e��w���d�Q�
�; \e�ږ�9�f����)t�pw���ٽ�*p�#;ɛĲ��p&���r�+&8EJϚ��$;<�X,c���s؟ ��t>W�F���ԋ�e&%,���a��Ę=�9ǻ�Ѐ�*��'���hx�9���7c��A6�3��_�  �F�*�������@2���9�J�
T��W."����)�4`����$��}�~�/���Z	�������a���r�j6�f�^�z��V\���"��K�F��"}�k\��ٺ2�]�i����J���ES��?k�儡�HĞ���o��F��x{�0���.[�������6�}i�� �U�V~.��
������>�^a�n�Z�z����,B2��G�LW�H���}��k�?�IAl�z,��gk������I#w�~��������g�R�� Ω��{�q�J6Z(��mU�vR��2%��T�\�wE������/��Q�V��eՈ�u��a��.ҮdP;S��]��(�
)�����)�b�)��P���oGײ$��W�΄�5i�Z;���G�+��ۄ�3}���7�F��Lv�"���Va���;��9��*��ʫB�r��!�e@��ג���)#��6��HyQ������%��&��ˌ2ފm!� V�8y�2wG�}�2Ӭ9 Hw�E���$U�Z �^���>�>��b�+*p�J$��]�;�kx��[j3=�G$lqj���Q�V�Q��h.���m;
�'�)�;�c�ۻ���
�A̳�p�"%\�λo�11g��A�{D!�e�;��aȌS%ٻ������6�̻�>\�� ��%��A$��'�a4�]�Q̆� T�ӫ�)>D �L�'M�H�"@��0P�\W�f_�3��+�WZk�~������YG/�ϥX'&yo�A��']�Ӷ$�[�~�C�����݆"���⃍�c�F���k�X�'���6Q�9�����-�_�"����v�	h}�4�o⻉)ʂ�Ӎ�^LȦ�
Y��9v����
��gzm�Ǜ�*N����m��?��P�%H�fg���V�;��Ln���� �$��U��EP��G���Al��p�S�����R��ɭ>"�A>3����{���-�<�d�`��EՔ; 4V(w�;��w ����H����31 �MN��Vn7�Q~jUw����Ф���D y�����9f��7�����pZ�ԭ��\��m3�C��J�r;���*���z82�v�l�.�4Bu|�wX�X)���W�E}7�
|V���/�M��u�iz�NQ��T��U�SC!Z���#@}�iש8�A��ɏ,y�.��_WM���@�8�*����ֳZb���7��g�)�����J��H�؈X�F���LޜC�&,��W�3�\+�3t���?��t?��r(���m6�{%aa�]��gu�muՃ����s����I1�iˈ�Xa=�9	�Z���W�Z�o�{!�[g_޴���:[��]�4�.ȃj��랡p}���.ߣ����WC.4}A�J��II�_���uEԇ"K{��cl� K�7��-[���3�����;mS9	.cu�(?�w�7�+9��>do&��,��/l�p�ce�b���'2��2��՗�:��2l|g�<�	v�l���F� ���O��R��@.ߛ���ɦ����Oe�s�k[�D���7��X�E��z�v��5����Ro�IB�::��&�IW
��2�Z��l�hΔ����L�~�X��۝p�M�$GBj��
'�)s4�
`�Z�㆝��vO *���~@�K+�յ���u+��)�bႂC�/�30��;B]?lJ�u���F�;�?p�]��94�Zw�ZD3H����hG��T���)2/�X�#v�����>�,��r4�&'���#�jȠy�,(A� Y*���벨D����3z��^�Y����z(esAw�zV��:���1�<�g���!�qo�ӆ�L����GC@��"J������,�V�;�R��`��U\��0�����1���ǲsʀ�X5�*��5I\7�<m$���<�Tl�Sb��W7˺�=���/÷����Z8Ľzk��i���k���c�8�|�����&su�������;
b`.���FטH��E�(f*���D�+����0�RX��Dl͵
&.	������L~6��P-�(\��;�nY���.<�i_��8��[����ۚ�2 �$�t�"RF۷4L�	ލ8[G(�6}�����ud*�:&��1\ �JA0ϴ��x�#��)�A��{#;�f��\K��l5�������h�:`��V��S�j�S��pĄ�����Y�6��c�>;�.8�J�㗜������ZAM�"���UA��l5���'�n=Zɞ��V�$���(��1�ᓛ[�ܰ����G�������f(Y���(��i�hL�M'Ox����Қ��\,+�#�ϲLGS0�o���8K� i2���9(�F��Y!�UV��I�>��_��/���>�[��y&v��K|�Z�\=z��!���0 �U���,$�"n�ϴ���j0�'9�j!���}��~�dE���bb^�A�:�.���WMz�h�)E�mi(�'��J����j�w�>��P@�"VZ�x_�ٓβ4$W?�A' O�Q�'
�aqݬ&v�p�.���3Bhz�*����ӓG1,~�iH�b��"ҫ�}��� ��8�O�e=G�9"bYw���1 oӿ**����j�z���!ӎZ����Dz�8a|N*g�OZ�R�UA�d�V ��?��]�m�4���7RҊ������� �x;E�*��b�OF��\�r�eae��Ld�����*@Z䄏�(��m[8�	� ƍ�ҕ +��sQ��(�s�-���"��Q'ol!8ĭ���_�m��K�>�
��-rt$0���"GǠo���C�1Y�.�����޳.�ԃgX"D�p�v��>��q�3�7�"4��:k����f��>:��aYզw�����I٘T��
5�ψܭ�������j�c�_�,V���v�l� >��j`�Sk6s��J�:Y�ڸ0���b�-�H�KØg�Y��f�Rf٠y����77U�J�9���sV��G9܇p�7��3;T������td�a�-{��`��E��J��\OI�u3�����`a��;F�9�E.V�.��� $j�KV�*���ą ��Q�?N�g��{���i��V�Q��!3�v�?���1��