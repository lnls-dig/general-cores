XlxV64EB    3227     cf0љ����t>Z��׭2�z��=�,�A/�A�*O���{f��v�����hC*��ҜC����� �?H7*/�8�4^P�O�K�N�@�G��V[�{��	y�Ǩ��(SЀ�ӛ���3}O�Zw#�ˀ�&lN��	O�l���1p=FD����ً$EҪ(���el���ᝒ�,oɝ.Vj؆������Rxo��	Qg���� B� �D�?d������y3�+h��弘��:r����Q2
֧XW�Z/�ҫ�S�\ĥ�M�"/��#�.%�7�������O8�>�A�3	����=9i��~�J$z����`w�gz�����c/7��d� m��=v(|�	���&1�@ν;�??P�T.��d,�XR��_��3O3'#��t�E��]���=���Kvwo��r���<�W�s�Q�/���/� �7��hZin1�ewh	x�rTEh,lM�v���A�U`5��g�Z �Ԛ��}mx�ad(#%圣����r=c
�l\�n�݊3SF��8�j�Y���coE�!�| �9>�g���\g)I\�(JYX�qsH��<���������K�e��LQ��k�DkB����Нȳ����_;�|� MAW�V�.�lV�0b��/�bEw��!����&Lw� ��O�}E�,z)��h�W��d�|���X�Bq��W@:LU<ǋ6=[��j�|�d�.~N�җ�t���Y���%JC�#����K�Z6d+� ��	���]1^��f.�=x�4S��3C]V\���� �+�����V�o
��Y(��������q�4�~R�R]`��2�p��9��/����H�m��D���c���AB&G��{0��ψ��i��w)"BF�cZ��t �m�� ~��2�W�m��/�%�gࡡ�h��k��ⳏx�JO,�S+
��?�Ȣ��Z%M�qxtbb����I9�z�
;l"���Iy�d)>�J�#��mć�u�1%l�Kau���2�a���m_�k�fp �f��I��Xg𤋮�s�2�6wu�|����L�R��|��*���?��?�ֳ�$=N4R���.���[)��o���s;�=*�l�ϗlp0O�	�Q�9f�B��{���%�����?�T�{����Gc6*~B�J+��tQF4�E�Wk�O�D��: �^�b�xl�ּ�8�e��%�ŷ��H&��[;3 �SF��=ܪ ^�ILMHg\�t�Fw���b������ �1E�#!w��1�F��>*F�^,���"�:�+�Sx`�s�]n��z �
I��Q��G|Y�涌�>j���,}�.Ҭ�M�����M�'��b\K�N�&g��G���M{ӌO�tb
%z���B2�����Tڠw��5qV�Dm0��`�9�s�p/�x?,'p����W���ˣ�Ǵ�$�Q�ML���f�/Ha;�s�6s��7w�,�q��d<��=O�_�A�Q��ip����	*CHP�����~��Ȧ}�ʗ�p43�5]�����VxD��=R����T.ݯ��T����uI	����4��FZ��{�~bN�V�c��q֛�8w�ڠ�L�P�ނ��b?�F3�@�K�Vq�1���?V�Ѣ}��]���ei���C��w��j	A1�9a�ҾiE�KR�O�W��U�9 �]��̺�i����a�����r5�Ť{/�N����K�6  �&��;��'{�Đ�NӁ�7�`��T��&0FV�ٻ3����e
����sn�6�Yð��4��4���uDZnj} ����@cD�A�-�	
'�/�騽��[.�q�5��慻Sr̅qzl�8Ψ\=7�a������W��Ţ�X����[p~4�@�&3F��N2x��&�p1
��3��.���iY'�򫷊H)G��q(�
DU��!���2pF7I��p�b�0��NԵ�������A�;�F/����j��U
U��r\�u���<�"���E@}��]�����#E�����TB8�rJp�.�)��|����u���\�n���g��!-z!-����]��qޕ_Ko��Ɉ�=-R嚰[=V,���w+��1�x[���_|�'~r�^>��搝TߢT��9ø���S�V��p�q�C4
��f�ι�iv�Y���9�# ���he,R;���h�������}�n8'���ģ"R�(z ��M�Zi-OZ8�]
��O�V�o�S��,�ݽ?��x�"��$�Q���w�/s�{��[����.nU�zt���1���W���eQ�P;[�9� ��?t�9���*���~6x%��+�Q�bў��?\6/~xcݨ�l������|�62�������Wm͹n�:l>���颤�8K�~
qL��tHpj��+-VϜg���;Q8����������'�e{���vcu?F�EUW�̛� ����JתJD��O�y���sN��k�d�؛�A���qa�MR����RSmRnN���Cs�MF��x�DW�At�9G����T�E�+D�=*��KA%���J��3�XJ��v @��D��a�I�fu%�'ԓ��$+w;l��������}��}#</�@8-��Iu�+�q^��܍E\X��o��i�0��zkz����Y�q�Sw���8;r"=�h�|��o��;.�[D���Q���>)�R1��iF��YLk?*�yg�-k���L���cAܠ�E[�u���Aј+y�p�Dڏ����,�Q���,�0#��v������7P�$,�NO܊ƭAO�k9�۹'1����w~":�UCݹ �sQ���d���M���e�������:�M�6���]���e�=e$~�l��v8@M��RmC]�G2<'��}�\�r3�-���� �쒁Я�-V���}Ժ�j�����I:�<�`2�^K�(֪�[Ad�����Y�:|�oð�a��R|�"�s�X��>��h5��^��+��za����8 ���N�]�W�ET�H�Uͻ�i�a՞�W�T}Q(�\��f����Ec �� qa���H?������yš��A��N�)��h V�w�c.^�P_�S8��h�gEOG���֧��'ǐ^��)�K��@z�����C>�D~���/�'ؤ�ǜZyV1�]UTU�-l�EÆ�C���,Џ[Y���'��v?��� }�����;��e��^4x?���,6M��S@�F�+T���Am�uK�h�
�N�̜d-+����H��Hzk����Ue