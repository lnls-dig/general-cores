XlxV64EB    331a     cd0��Z���ँ6��D�9�)/���G$����4�+�$�;0˘�z�`{�S{��K��LU�&�<8���95���|Y+���D�ߧ�;�1'c��"��O�9"�����a�4�/d��o�>Z7�v%��������G��+JKZ�)�;��Z�H�Zo���{���벟�И�yqy	�����yMKZI��C������3�Ƅ�:D\0��C�#�mz�*-c����U���F=0��vFc0��Ʃ ��)�5mx�zO-��@?�呃d(Q5lT��Zf�$Mfnb�T��-��gi`�,P�N�TF$�B-ʝY�|�E�'�q8Qϔ��R��~��_�@�i�"4K�i�.e|�=�����+�z�[g�u���|"�Zr0^ً�.1@B��ju�G	�:d�@�P�.Yf���3H���!ƣ��'�1Тa��,j@-�cҵ�|����1l�Y_� ��c�Q̿�lnv����lǗ%��ZC�_�6{ǐ��֙JQ8!�{-��Q��X�Q.����i�:|�A���d`\��:Ie��rn�����wc1(���3Aq+��j��iE'�z� ��o�w4�5rՆRB�Ix�5k��/�6�y�M�>Q��ǋ����hN�#:��iMp�f��$y�>Fm_8�_N���A^%J�e@!޿��~��fJ�YfL�&X�R�!���*K��i>�k�EhD���#9�/6z�y���/���X@(�UAt(�'���,i0*-�v�a���n0N�C�?]!ȴf�_B�,K[�z+_0�J(���A4�N���Z��%��+�P��c^3���y����d�)�"�P�V=�� y��$�%Ʋ����2���6`���w�@����kU���6�s}���8�.�S5Q!��3�{��ԍvAaEH��!G�J����TV��*n��4��r��l��f'�F!�5^(�ʌ?�uK�A(�c��-#��c�34�}�jJ==k}�u��]�1t�I7��������l��Eq�@)<B(�Tum�g���>��w�l���j��'s��dcs��R,
cg�E����6�?d��B#��2!8*yK��)�����:������`�1�d��U��9
i#0����{$�7���eW^����6�Oy���3:o�ܬX���S.������,�i�;Wf�Uc��X����x�$ �[Vc~�j��n1�̅��>V�y��'m5.�{�6o�I5 Lf�~�h	�Uہ�O��X@ΦA��� �b�YkLRq�s�YMm�F�|�X�	O���1>�</ �B���gI?�:��I��#06V�>��B����v���.U�Ѵ�|� R�����������h��-m
9�K(<[����^ߣ����1z��j%"-�����6Y�J��^f��+=zL��-�>k5�>�Qn	9IJ�E.Iu˧���R�9�6R�����X��N��SG�_򶰴�Lt��MF���q���<�J=��a�H��}�Ӭ���f^��م���0�W�veM�D��gm[���i�Rد��=��N�+�k�9�������.<�	k��ݩRǐ��Gc�µS��������	�1��1>b�2^_��bcg�e�&Iy�r�y�rB�\�y�j�U5�	�K{6yՖR���{�:<!L`�PNΥS�U���;	ҜՈ#	!�hl(�9S�}����4�mz�GGwd����A)5�/`��_�����+�P��;��o�l[���)�(����� ��*�0����|s�����!WͲ�5�첅8 :@�-�̬Oǯ�!M�޵��3q$-�����5$#s�d!�=+��P��mn{��:�`��?�L`�iCkVm�@|z��A7/� }<�]V��u6�w�F��|��$�伷5��> �����T$��;�E z��٧�1qJ5�u�����W74Dy2�?��I��5!�>�������>I��(�0���MLJ#	C;O��wb��o��W�iI׀C� ����+��~���oR�	�^�@&�L���g3+���o�4�vkяA�|/߂=���0���jq�T�,�)��s�5��𓆃���	"�������(b�"�-\Ӈ��P���T�q������a�A�6A�LNYg�4�[��)�f;uӧ�q�F@f��ÈG�:`�YB~�xD�Z��Bl�'��h��r�Κs2����g�������z���)p4x���=�aN@��`�bp�	?��I�%Vߜ�9Ҿ[������箙�:f��k���eԏ�57+�mpy����j�z��k}�̢e��8�����J�>|
�BA$���?��5ʩ.��s6xI��	Y8�K?�b. .� �?ٌ��*�\���![IY����㭷�$��%�=6(?�럆��0Wp�%a�Q��k��J}�4P*ߣв}����ʼ��!G\p�me��oS��!@~�=��=��<P��L�/7%�+qTg����>fX(�T|�}���u62��v7zYp��<t�W��|�&l�^Rߣ��GR�|i��ϒPn����X��)���On��J9��H�����O�L����6F�&^[�Fk��� 7��O��R��ؒ�q�{ӓĵ-
PG��`�kL�(���M!���]@�-�`�:�J��F]�=�jN�,ST��-��+8��߰���v	�^�i��z��Д�tZ�Y(ڛ� �����Hd�h}�2�>Cȁ{:F�Y���ѻ��4���E�5,�-��]O�V\Q2���)�v�Lbf�r7m��1��`xe~���_�X1�aC#
���t-���XO?�	m�3�%� G��%�������w T� 4~��>�y�̂�|���0��2�Ҷgg�J���|��RJ�
�iJ+��A��k�y�IJ۴d@C��B�����7�F���W��	MC]�Ʉ���iB���5T�{z�w�+��(L� ";� �ԲzRtMq���z��"�������o�g'��qC8:-_:��%4/�W��])�9�2ɷ��0&G�Y�<�Đ�����y,eQe�Pae�<]��E�ڷ�T=����b)e#��zv9{�[��vs�Z��%����â(�-`g��Ȼ�V���楝�0=
���ݱ�%&;����u6���2z����I%�k�m�q�u��Ϲ��������b]��2|b�֩���&?