XlxV64EB    c90e    1e80��X��i�޲�ѵ�s��ؐ�|�5�x�C����;I�x�W�A[���c�Ōi"\$���������%��Y��IH���/x�̄3�d�x�rI����A�r�l��A�i����6�q
�Tʹ �G��rR��ps6 ��/E�3�C|�s�E�X�@�ew!=�H����T>�Z��R���_�q�$����i����䓛�J��G�e���X�x�2k�
���iT���+UU]??UJ��pL��d��q=.������>l��B̌���\n�
�X�Jy�= 	��PO偫1��!�Ý�m�u ś�QQ@�V�E<tN�����?U����O���H�ѹ��N8�u �|Q���dҐ�����J@��2�ݻYz���	x]3Bpcs�l����M)9_9m�5.E�4ٸB����LG���E��At4	�7��ώ���ϲP��.�n��9m�Aa��3�����	ؗ�MZ���6�@l��%�?�Y�V�C�W�0����H��s$�����ݱ��˫�Ҟ���~BFG'�N�>dY����r���X��Z��lU���l"J"�n��D�Sq*�N�x?����;��u/1Qm�EK��fI��c�H���;�@)(�-iw"^����ɺ����~�Х��s�V@��D��y�6�Lp��K�e]���/��vL?�I����|����8z�� ���h:7��V��F��>'�q��Bɺ��	�n�y$�w��ͩ��	��Rla����ޢ��0l;#��_�n���,��黼���k��i��GmME�X� T��z��.����څ
7}66]"���>��O��q^g!֐
B|B l������[���fO��Y���ĥ���Y�
c�B+��׫~	{���i����H��58s}O.�s�7�X�7K�)r5��>V��,��Hc��YMu+j�
Q��$"��P�(��Ja[�xM�pD��1����~)j͘7��6"E�n�ԇo֌��s���H�H������� tXA��,�����w8��g�gR�s 4��+8r T0�B����C]H���$��������dJh���/���Htfy�$ٰ�� f4�IH��E�9�?�_S �\Ƕ,3ѵ�d�9��~�"�,�)�0�N��~ջn
�Y�)�����w~�^��4
�`�}����,5�����B�@��M���5x."l��� ��.;_$�f �BFn{��QWA�3-�a�6x�̈
0~���," ��͜2���Ap���s)#��N��Z|$:�L=����b毂�
^�>��`)~_�^����l���w��B_��J�pQ8��[g���϶ċ{B/�w�'zl����0�x�0�zEQ�c  7ŁH<o.�;�(~%O��h���1��hO�3��%�x>3B�������g�J�|w��!n�h�?��ClҐ�b��C���Y�=Ne\	��0�SXG��H{ @�v�o�c�؀&
�Y�Tm��9����J
t������+���V�4�Wvm��W��5d	�!���*�y��-c�]N�[p?3��G�{�#���m}P�y��`g,ku=�̓Pj8�4=�h	\��6._�뻳�Ma(K�>&Do[����<ˤ#����E&���/�5�x.6s�8:�dSB!r��6�i�brt��X�@����F��s��4}l����0^��zP �!d�*��7^-�<��j���%�*��{<�JxӸ���
�u�kD6ݔ�$�'K<�6fE"��5g�p k�3$
�]�,�k9�s�|f.���{��L�5�vu��`�% �M��Y�]:��4�4�1�UQ��05X�_��Mw�{a���wM���e1W��H�����<Zl�?��Z���E�<"��v�.��W|���*���R�&��v<���՜0�Σ9G����m�WM�~oxH�گ��etR�n%c���z����[Ηj�CAh)���e�*!5�'3�@[Udg0��Z�g�&�ax��Gfss��e,� ���j�	=�1f�Qw��m�X>8IǔR��t5P�_@�������tskDz̃Oc�m0��o���׈�Ʈ��(X c@6���h��I�D�"�� ���vhh�b�&{������ ��+��,L������1��UIܮ��бcWj��͍�fS&xK�,�!:�R�@	����,�ޫ�)A�Urj�z.���[�j�1!@O�6g�_+���R�/~#cT�W7��t�g����\	�P������7��[v:�`�D���B�i�%�]���^]�ECCg�������i�& �׭J7߀E��C���b�;*������g��o��gM�Y~:/㢯H���Cڛ��.� ��.�Ӏ:��9���;�"��/z�U���O^ʉ��s�s^V��8�SW�wH�h��7w�M�'��!Zl��(�9�o�pYp�!� �>����0v�Wkf�>a��M:����������{��#���c�L��7,%m��h�i�FE�������b��;�2��'DkZ����\j�d�ɮ[u���1<=��dꥅ~�ս"�mu��S��ϼ��DE�e�5F�}�7�͑F^Q��!A���w��B��A�!�_zO���U�Sä1h�,��8��Wiۇ�%�֘5���pB���9����տCO}C�F����gO��Ar�0C�������π���D�s?Z4��,��x��!u[�7��0;���i$�����Z�L��y�`�o�����ٮ���}�	����Y�g�T�𤌯������|PO��=M�YtO�Lح,���@��|
�2����j8.W�t/����w��p���a�{�=ܛU�3B��&B���V�0��z��n���l����߇�B�KEg�#�(��~26�O�n�EH|��_��"�]�e]�Ա��s2��oM-"lLeS��AGӑ�f?8������@���ʦ�)M���^�������Q���a���s��u}²�p�������!��h����K|nI�f�Ȋ]G܊���P0F��0���h�󪝋�e߮�m�[�1Wz*>.��_6�y	uԻVxl��8i�<�)�v\jԤn���	ky�a
�� �g�59��5��
���0��f��J$-d�����/������nr��,���R�*���-����\5�yS��$^0]�(\��n3�������o�E\F�znzu��S� -��1E��D�;%�t�4�%�f�'ւ>�� M��MBl���@���Qq�h�)�~��IY�o?��틙/h�ڟ���,��:�	��UWG��uX��!�-�'�S0����� #�J�ZN$n;�\����{"�X2i2[7R�
�w٣���G8
���b��pd�S�)m"��Jд���8����+��`�{�%l�ۜhZߎ�͞�mV�y�B<7k{��K������j�A:�2`'�ǚ9������y3/@��lFo�z7z�� ���᫄0������"	�M��(�>¨����@ޥ�s�[��f�R����]�������ۉ���c��̓�;�'��|T�-q�k��n�KLU��@f?��H��+���:;<<'"�DG($A��J���6|�� NYa��o����E��jMM�
Ib0�O��--Ds����ˆ�y��J����GK�6���W'Q�`VO��$͎�M�q��_�St��K̴�`�9 {mY�crz����@.!Xo޸h��=�[`�ᇁ�R��A}s2R2���!��<]�����%�7&l{'}u�o��8��}_����*���lti��@@�o-H����[{�C��t<�%�/"���\�����2���*��\Зe��7"	∭6�H&��c�:�;��I���p�Fl!��F�bbw�U"�G�A�F�L��ū�uy��Z�� KCp�c����ރ��!�9aJ��E��>f(��Ш�9����P����R�??c�M�p�{�f�s0�3�G���u���G�6z,�v̭����FYC�3g�m�^-�E!��;���7��t�?QY49�?��1y�J/D*cQ�1>*\�y\�؉t&~JƟ��<����j�Z��T��!�=�^��N�f��ޅ��H���k�1�]�����}~�Am��"E���h�/����([޿�FGt}�i�޾�oGҭ�~�@��`C==�lQI��������Vj&r<��&���dz�_L)Gm��Y?�cL��$�N�V��{<0��P��.;��,_}�x�=����O�ȩ�lo-/��`��E)2�򾀅>e~ia%�|� �z#H������b�I�߁?�No����Yb{��}�0�R5�K4��*��g��E-��)� ���(�EmR	D���6u������|�i�G�yӠ��-v�1{�Ynv��E�ka�Y �E\Nf>g��¼PP S�N�vC�{�����^t�G5���'��a��6���´r��'�=΢Q?�s�k�$[c���O/��u��D�_!�/��4��]��px�e/�a0��8W֨&�1d�V_$�/� �"$	��@�lJn�)e���ʰ��UZ~��)�}z��|��&�|�i����i#6� K���[%�ᎉ��Н�ɰC1Eɦ@��`?��9���_;k����G9dk��E�d*Ja��@�V�����4yn��q��]�����o���'��q��8/���l��g�"�J�O�su �9���l��X{�x��-��S�&�#]�J�6(�z���f���gǷ����U2���Ps/�ESk�����d9IC�,��|�{
c�@�5��J�`�<��Y��5?�b9W���[� A[���_s�sj�� $����_�����.P��v0,�#�֑uy��;Ȳ��D� ��~X�Q��׋ڊ�s�|Y�[v�'7��̡B�?�GM����@���O�
MJ��gddiiq�5�i�	V��jњ��c���⭶d� �d��DQ3/ax?� �AW4�`�Tπ���"��*y��Y�I�{��j�S�p����*s���L[l��T��SL�mnt$[�^�S�iut�8��}��e-�Eu�So�U����E�a-u�-�Il�w.�j������T�⭇�ĺw�6@���l@c���y�2`�yQ�F�C��	z�H��� ����E��'�@1N�, j�
4?�O����>w��b���F6v*��n���G9�s#��Ҷ�dfDp�P�&��uW�����Tot�4�B�	��8g�.� ���`ƫޘ�+P�f�ΊTX��EM���r�!� �p4#�j����̝��_�c\�F�l�����~�&wѠ ����cˢ�[�c8vS�� ���{��$����[?)$��Sf�����z��	�������s|n����AR�cgtB�v�U�佟�j�d�^�v=:�
�����U��[s�e�0C�����8D�.��=<2�Ȣv�.�ݍW�n�޺q-C�Ll�U`�7�IO�Eî����*�S��G�m-�����v��^��N�60n������`:�yGL|HP�Ȭ<����޾�]�2Fn�O\�80�f+���y�B�y�r��z~�q\�b:��p�£�>��;p� =��5�f�'�-!�-��J��DAekn8��\�d��xC�_�(��r��>����v�0�ך�;:��Y�������\���}��� �yCn��⿉��͜g�(������GOb���/
j��{���i�]���1J%��{`�lք�`A�<W-�O��U��ą���%R�=]�W��	~?�d@�
VtEǨ��߈Z�ޢ2D}�[/tG�px�ȅ��|����Oy�\��U��z�d�����CZpRZ)��t�x���̚k\}HaY=�F�2�%I׎�&`�C��6G�ut|s�p�D�)���-j6��锷i�W��w�����s��W�U�A;tbIF+L�S�HN��2��xx��E��q�N;+7�4@n?𥉇��4�l|&6�4ܲ)��y��6�Y�W�r�e]�o��1�k=�9�G7�'���I���X�	y+�P���T�÷L�ϲ��0��$-�ȋh���@��<����@�{���B�9��&C?�', T��:���|�hPl�7�Yis�=]6�{B�!�X���i��A}]P[������f�&}U���e䈗8�>=ЛT;O	~5k��.��Sz��(���5ډ�0��
�*�ﾮ����<�
�a�Ai������{�`�A��a�%��c޼޷&�ߤ8YI_��W�f�t���U��I�"j2s9&�Н��7|���r�7ƞ�d���%������r��Cpo�D�|T��,��j�C��c�@��9�M�ߓd;��s�"���&Yt��RR�5�,|�Ym_'����c> �Z\;��J�:^�v�-aV��<�$b]���FH��O3� �IKo���xiq�)Ï>�Yn�ªo�j8=KM��O�20�����<G����#�]<m�a�8}���9�ԥFy�p��
͟'��v���	�:�B�/�w�B���-r�r�MZ��x�?�aV�1���1	��z���YFR��%w�I����Ӥp$7���
W�;0L��V������%[�6]b�|+-M�����[a�d3�B�����ق���"�J��D5��捕��}��Py�.Kb�-_�'}�:TJ��Bp�	�NdF�����u{��� �
�R���P
F��֮��w�y�ogyZE�B��yߤ�D�-eL��+�S��)�͟��Qi<D�v�C�,w�G��wc���3�j~��y��rߪ�oS���eO*�(E�QX��
T�(g��N��6I ���G;�Ư,�QN�{��&�X���І�l�?j1\������������4z�f.j:r��{+k�kӬ�����rt=��e'.�g�y)^�A����#H �}^��b�-�P!�����s��A��6��T��)� 5�x�a�RR��Gb�mZ����w����0^X�V/�ѭB�`S��*��0x8�;-A	�Ϛ���,�a/v1�IC3Ș��i4��&��1��P#��$M?T�9�1�BT4��|y؁_�8c���d���{�2hbo��\i� 0l�b��tU}ԡ��E�顺��V�xrf��d8���h���%V��� ���4�8<�>}��8�����^R�A1�i���~[w*c�?b�R-�H�6�XK�Q��5���:F��z��ر�)�7��c���2c5��J$�Q��[�ʱ���bt6����֊���z�t�\ ��k�W?�.���a9� �Yz
N�������DHI�2S��(��&e��y��OdXPp�e�=e����\'*��pCvӈ���C?V2���N���K�j��'��=D�V
b�>LdU{�˃(�����4����8��[\�B�yu�,ё�`�Sоh�|j9h��t��Ɏ���@�_R>=�aA���D��d�1���y�ca9�� %�R�Z�̼d��z�	�9P��h� w�pQ[a-v���n�my���Q�v��n���&�w/�9�w;�(�8� -{ID�m[
"�` BY}.�������w^	ډ�����"�»��n��É���rs /�5W37�4�If \���Ju�Y|"�g͑���@FS���)���Tv�]ށI���0<4�}��