XlxV64EB    82d3    1750KM��|��t����$������鵍�uZڭ����Slt7���^�BȎ�3I�F�y|�#3-o��D@�%�5��઱nWfĕ��~.x����N��Q�j�n�wǻ�@~�m���ͅ��P9��;2���ư\�E��mo�iP읥᯶��2Q9�j�3a�(	�Gmʧ�n6�§�<E�2��(���i䝄�#����;�BeI.W3�|qֆ3�y������V֛mظZ]�o˔:q�e��I.	�}��?(w�\�U:�����չ��/�jw����w�"��!a� ��r��Nv�2F��?TP�f�C�n:�W�Uφ8����y�z�vV�-yv���l۳S�t�W;)�J:�����X�U�3Y{ɍ�ߔw�S���oF��aSy1H���t[����@+31��}z��,�x(��}c�p�����n���'��~3�@'��K�%��T�R��/�e��S��$ï�"��z;������k�L���c��v\�-&-�3��qN���7�z:�Y�֚ha�K���B�����O�����/M$��=��X2��m�Ɵ���������rCќ�b����{�'��e�ٿOt�@�o���v���[+@(Y�n@Y��k�}^ջ��j̡��_ȿ����o9�B�K`���+ÑI_⠣f��*v�Wy���zӘ�B������,f�=#�Q8�Dݱ۳U�ڔx�py�_�:2���♜qNŗ��K}s\�$���sb} �ƪ.��
�6�@�K�1_���abנ�N$�B�Ӭ4�G��F�5��6��I����%t�d&)]:_��1@���<�aX=wk	Q*��B������T+P�S����=n�"[�������1���������n�Iȏ����p��āLMf|��l��@Ȁ�{-��_-�V�!��p��,;w)��Υ[�![�7c|(U<��ZDUH%�8��IyK�q��wZk����4�<�����?�����wXl+-�5��`�y �+k�o
K�\��>O^2<�v �RW�r�n��U�}��K[����^ծ���Clv�@�Xvw�K!�o����Q]q{2�u���nI�ʙ|V~��8*DN�#6���E6dp���T�����:� R�b��8���4^p@2������?κ��%Y�h��<ø
PVhm�!$]�x'�Y؏O���/�v1���coS2�;�0�q���G�z܃�ӵl�O��3����2���p؇i:�� �6s�G���8�x����P
 �-p�͝�AB~��3��ݽ9�h�(p<U9*N�F��D�Z��W���ʑ��8�dT��;���HP@7�`���.���q
s�˂"�g����c��8�!���5)(��7i�ə,��"a(NS?jVz\T6��=�//�~�v�	F�$&XE�_����2�lT�%�C)`Ly��IE���B��K;�lIA�L*�#��1� ��*���hEn��t����L���j�P�9���Ч��5`�ʢ7J`��./R?3by�5Y���{�XLi�7$g�Y󥤤;����.������vh�٢��Ȍ��֝ Or�A��+F�K�u�:�p�����a���[91諀{sߠ���h�*P8 |G��������U�w4��v�ܭڸ�O�#���"�2hq�K�c�����l���yMK�vc!����j(Y[I�NǢv�&�(�`���8�%Eʐhh�&CR�0y� g����~p�tW� yM��Dh\;Rnh��<��/�f+G��Ҍت��cS�q����-����(������M0��u�*/��F�"m�B�������	70��p�WhvC`�?V�5����.,�T�����YE~̶rUo�j�(�4�����tQ��[Br��u����͆����о��6�z�@e��{N��6���0���D��$����*�F�bƃf��T#����Uq��&/�Z�
�K�ه�^�����`�<���3(x�h�vZ�"p���1�;t�cK#��Zx	��>$��0X��\�aLE�*J&��k���m�)� ��D�Ñ�^a�J�(<H��%��)1�����vQ�Jo�u$���V��W YYM���ͱ�k5yʩ�ך.���~�x/\�|��ޠ1I̖��,bw�gEq �#��� �⨊�hK��yA���y_5�=�&�ݪ2��}+V��3(��>
9�}��[`%�R���ʠ�EG\�9��f`:iK�"��Vl���S������H�ĳ~ �/�G�^0�4�q^�"a�b�ۦevx|~��^����PO9'Oۗ�1m�b����0�K0_ �νfk0�[lV.�8���/���
d%��_�"L/��4{�'���f���"��D�����gYm��,o�z��9���̅sV&�O�K�_���`��a���%T�b��5h�$����f����$�S��YR_^���8���'�m�e�0�yr��]��``M�W�����y�zy]��\O�b3����>9
l�$b��ł�
g�g��h��U�}d\(/��+�*���A��m�Q�-�g����>�׸9l�|x���.[�ܧѳԊG�HY��؇�v[�\�&l:�L���lV{`y���E�xjÆ��
(z�:�t��T	��>g+4��Z�2� m��n��#����M*���/��_j��h�toX-������hį�C1��&��~����NW!��ލ<:�� R��s<�v������[oz�I�ù�~��@�t�:Xb=ь�eY9(�/AH[,�kq2�mFhO�W���r<���Kx?U�]"�,M�R�0�7��n`���D�1���@��jԟ^Y`�8�/ƺ`M]|��BNa�Mh�y���ɜ���s0%**�"	��.��31X�X�!��27�M�̃V`�q�����h|�aS`$u �#t�8E@�귕ܹo�JIQ�2\h�>�|�%HM����-�1�|T��zK/�9][t�� �P�1I�ܓ��p7@p��w�� V�
���N굫F��c��u�K��4E�Q����� I����T���:�7qή�7"�� ����{_)tbM��\J�L�o�?�Y#� �l����Xy'�s>�*����N�r�b�M�0ػ=ѷ_��A�����'vԜ���F+�W�� �<����%��1��{�r0�#F9�VD`�cs�8�M�{�z����.u*��To�Y�S@�#D\s�8�#�;�IZJ�w�͊�{�[�&<)�5��v�Ƈ���0���?k�8�#���MN[�'k��s~�9 �<�k���b=�/?�ҥ���3����!��<�� �z��Wֆ�l���J�I5Kf�)��!������_�h�9
�$߸v��h�ctTM,���g���t��
��?L�N���o��}�H�����y�j�n�~	�Q*�5���eRן&t����0猄�o��`�p�,�oz����(�<�(U��K�IÐ
hc�\��M�b�������
�B٥�6�V�Ir����p��YvC�]LQ�7m.��:�h��������A���+�fÂ�Ox(F��x�L`߀��g�7�I�0aޓ����ŕ��p9%	'�3;��F�A4�(�/Ɗ�R�G��`�$#k'���e���hH��!{�.v�w�i���n�+��.�ހ�2�z�'ëpki�\ϓ"^��l�lB��t��F@��,��Ő�dmʡ�����4��9�5�h&K���V?j��f½��n�x�ڮ?�cwCM���!�A�1��ޒ���2J��<�U��3{LP�S�|^$[xWX���M6����µw�F|�^*����U��
�I��hq�)��Ni�_ia	p��k%A�%���a�r�aw��s2G��]Mh4�>���}�(�.�j���	I(-�yg�s[��,mC9$@�fr]��A��C��|6�;?��߲�`��J���43��<��ڔX��Y����i0���'���)�!�w#,}m%�؇��X!��z��7��o��zOe��UdU8��sO�-R叕k�:͡�`SO�����+��jQMUH�Kو�x���t}2�녀��'W�]�� '{FM���A}񓶦ъ�N��	#!��z�?�8�f�>g�-�F�?'���~+ l��ذi�Vb��!�Ε=� ��z���Av������}��H����WS)� (B��}41Z�E%�6˥�5�I@��ْȦM͊>�Ե)I��+�N��0���|�8]1I��Q�vI����w�?.#W�C;顬t�r!$6���'����ր`��D�1�|;1|�Ӿ�\Q2�������/�v��p1���9�����SdQ_��,�^��S���ݠ�e0`��Զ)��k���LH����m���f��x'�;(��/�z�B��9��5^%��cq/�FƳ�9�h��C���4C������<���:-Nn��2�E�{��#������+�U���{�e��4��x�-aҠ�^�|\�wu�^z��֯�����U#heO�b�[���ot����(;��J��ʏE��2^�>r� ���q�f�E}Ft�1�z�c�8����e��ȇ���o�k��OpB]WO[͖�Ж� ��c�ep�+$fv�T����j�I���4v-���@�H.L���1�1R�`Q������Cv�����E�&�J��a��-��ne"�.R�Tڠ����y��+6!�K�i�%��?^�3|?P�d���v�(6�rN�S��4�fl�&2�����"�]�9�m��<�dt�.R	�5�,3����:���򹗎j�0K=��$�_����:����ңZ�.��X��!V�kF��~`�;����(hK�-���o�:�M����fFo���?��K@����Z#��|�0�J���d��쨘Y����I|����g3:�G��f2�@,��w4s��Q�7p�3ϥl8�~?lh�~U�������C�^k����/�xӥ>�u�LI	��~��at̂��ղ����N��=�����ڠ�$o��m��Q����GVPe�'����*�Fӄ	��4s��������E���9ݟ�e�L'�Qpi�~�Y�PS#�˫���_��B��OZ��@ߴ�]#d�ҧ��|z��.��,�T�ń��;m�=�!#E 䐾�p5�Y���),q�*S����u�<%H>�3<�8"��F�7�H���o��l��$y�?���N@�7p�ɒ�a�o���`���n�����y7a0�&�滑�h��`q��"W���C.m���St��5^��פ��&�B�i�̤��M�z��i�"�d���A�,�P�$z7�|I��<���C�@�Q�7����8y1XʾN�>���1��N3$sEC*�W}��l;H�|K�ae��~������`Z�����P��~�)��;}����Ӫ.ݠ��Y��zJ�p�}�����Bɹ��e�lh�DxLi4#��@�R O���u6^��<��	m�u~"́��ڥ?A�.����}�Z����utx:��f�(��uc���2�Ȥ��:x ʹʼ�)W��fkl;�e���a���7o�l�"M����V�$�%�l6��l���1��.,� Ԡ���zea��r�ZFrO:�@K���Í�k��[0�_D$�	S�ޥ	6�a��);�;��^�����Pk����q�AWO���bJ�Fک�"�5B&eC�L�Tؕ�|�l�!=1�)��~�)-�-��"̿^�^P)g���u����6?C�,��{p�8U����o����L����7� l��mj4����PL�"6W��o�