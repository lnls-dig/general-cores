XlxV64EB    6c89    1840�7ا\i$|Q��<�{�_�5���7z�ҧߚ��N�&։!�sS��T���p��W'�@� `�3/+u�h�֧SWe�&'Z��2��L3y���̌e���L`�Q��E"T���]�����X٫�q�M��@���b;db�}w=S�6ʇ�V@� v��";���ͪ�}l�����tS����eD�6V|H�7w���f��(�ew��s#�V۷��\��o<�x�ڷ�\���/�	��-�D�q5�g^y��a����z�̱��)�ԌŲ8�(�1�K3Rĕ�L�J��7���_f~]݃�K3�X�V�o����3q7Qx��y��!1YC��z:��'�ꈑ�hF���ص�G�j�@�r����s��J_	%ޛ��m�I�t������R�a�a��v`�]J%�U���8ZƸ���U���
#�M��e�XY��>���ީ8Ƚ�䴢/_X��F��y¬�k���0J�����Z4,��¦%_㾏3��w�>=>d��Z8+9ۙ��I�����������t����㝓0ac?%$�'��W>Qxa�����U��d�F��S�Nm/��&������K�=^Cu��q����~��Q�d�;Q�i�A�L5^Z�A��e^�P�0�Xǖ�睊K��,+�t��`5੝zd��	w�D]:OP��\R�h1�tȓ��5\š�
�)A�L�8x��M����u)�nמ����`ܗ�Ν@�ǩ�v]3#L�
+K�������vs�$��u�������B�`(`[msU����E����"U��
38�?5}s�x��aԧťb92�~�.<���rG�+"��ْ)�>���3b�g9kD�!T�D����V*�i8��[v&d�Z����!@��gG�h���\��.ì�%�1̳���B4���ɰ�����X�U9~x���d�w��U.��=&��z��\��#e���Ƣ[���@�_%Y 
O�=Z�(��������m�s�N�i܊�F����!����"f�"1bk��x"�E�0�EL�uZ��q�񊩗P��Y��6�Y���B�D����+��J�GsC3����o7d�~�/ ���~��ۑ�Ǣ�t��ʡ�t_�"X���+Β�,�����kn�vO�Tg�����7R���2�i���G0Τ֩��sH+�ᘸ�ݥh���,�;��k�rv��&���Y��`��%3����]��]�v�����3;��f���*�^���a�A����]E�k��TgEA�7e+�V�U,A|#�C�-<�1E����"=���І�k�t� �Q��o^�_`�N�wg#�� ��f��{�Ҽ]C��>���^c8���Q�Ѵ��A��@�WQ���iG��99�I�pݿF���1@��ԥη�9�� ���L�E�?��{hX�:Q��Ղm5��scK�=O�}-$q�_�E��L���$R��E�I�M�<�Z��Ί��N���N�uR����>��Y�6u쇦z�-��@��&6��G��!��+��J��D�����H�/���D�e�wF�I�6�x _UI�p��5���J�:�RV8Q��z�YhT���Z}�@�0rT.�϶Da���ʋ�� P�4`�	��G�]��/�p�;�l����6����˱�D{��="1�vlXp��a�Z��b5�h[ ~��I8��v���~(��M�C���4N��<F�N˟.�s�,A�O�Zэ��L!�K����"��i��O���ш��r�!��59EM�+�$�b��(�5�L�L�+��"�1۩#�6��Ӡ*3��m�~e�*��Y����ev��D!�WT����3�PNÃF��a䖕M��B:�Vbi�u�O�Q][q�'h��
$v�0f��Yc���Ƀ[�}��_G�yc�.����M{*�@H�'fB&n�;� O'b�"5�J)�LS��~~�S�����D/Y�tI���+rzw��ݝ��J�G� l��N�m�E�ev(
����V�28����WU��P6X�2�����\����Mf��K��L�Y��Z���Z�6��;���Q^s��n/iO��,�±΂+�8�=#8�r|ޟO��΍�D�n���uٽ_qd�_>�5��9��Vp��K�D���@*آ�	A�,Zb<JZ�Y�����*���
��˃�i�ɲ~[4<�{�NB�f)�Hi@L�v�>M��M=rm-�y$���NU���6���~T�
dE"4�Y�����N��g%�c ��R�ʍ�U���Ԟ�p���D�v�۔��,��a�@�N0.�w1�*�q���ӱ�G�tK!�y76�L�;G��#~ʾ;2j���Z����[I�-�$��z���i&Bw}�'��Lce�b,���k24��U	�[�a�'��>��.zb4��_TQ�2�erbTӃr���-����-��j�J�S2_R�����O*`�͔"��};#8�瑶��ϳ���ls�Y��r��~t�Q��x�¹�l�0ꢷXWFA�@P|k�=5��p��x�ԿF������l�Tt�qU���_=�f��>WAD|2�:3����7�)(d�
�)�A,X{���=����"�[!sp�K�a��/�*��;va� ^�Y���N�P�ۅ�!�w�+�`���cQ�(86e���|#Z-�\f̾���z�(×V���9�V�صyIAp��t({z�0�s
w�B,b� �*
D�pMR�i���R]%���G6~��I `�ޢh,�8������^L]dCҬ3��Cg�\=՝{i�����A�pL�߈YB&�Pѓ̙	h��ݼ͊{1�7ఴ�J��,<AkLwe�=4D�2�g�q��y�.�Q%ރ��*w��.T��ڔ�n��B�}r���)]�h�M��ہ�U}�%���r_(YD1L�P���>(�Y[����+��Ș\��5?g_�6�=�X�ܸ��ޟ)LF��B��aEq����Nk@��y Z����ZS�,m6j�\��m���]N=�d��7�����w!U��������y�����i�l��@~��w��U{!O�5�K�Đ�f���م��R�jԸY�9�E�%Ɛ ��&�x���L�(Ļ�h��{���E��e'����_ܥH�b�����q(}wR������7җ����S�8�H���&,������%������B��=�����g%*>�A��셝�/�&g����6�7����G��v�[���!���2�_"�J�Z��M�>.�Q,M0-�N��.�ٞ14U�	��'�0��|K�{�Ŋ2�{ڹ���#���RW?�w�~�W4}�G��OF��I	�&c%e`�$���)%����ho��C���9������, V���(E�`�,b0��:��L;o۰�ub4Y�q�m��@¯��هJ�c��۶s�W���@���lHr֐s����Ȫ/aap6�O��;�(��J�'xIUC�1�o5tKL�qC\�&�*9���9�;���x[/���%�J̓�
0˗�ݾ�+�+�}X"��ݐ�g�Z���T���s�ߢ`�C�N��t�JJ����s;o�n�SU~M�>A���z�Ͱ�1L_�=�TmU�yKY�p�|���wЩT��P��TP�=��oA��V�Q���,,6?��NR����������U�ȷ_���&����Td�`T	�O !�,wA�آ�$�r9�)	���� 搶�j-<'I{{W����2���X�Ӄ���L
�.Ț!5'�Kr
�/��`�f]�x5�nJ���u[D�7���J�����Bd�x 5g��M�#���	�y��S3\D���g�����f������rX�t���ȏ���%�0d�/��e�?�Q��:Ԁ������<kY׶#�j�}f�Qb"���/hh����#��7�_��4����%|�4�<��/{�XyT��S�`o�,�?����1�+u	��ۃEB_���?q:!Q����}�P{�>�ȘF#aᜃ ѥﳮ��I�c�����3C�4�����1�Z2���^���<I�L��)?���sR�:�s��,0'�0tY�{�g�����-S�U�f���p���m�,����� Ѡ���]�oQ���i,#�$��eS�� =���y�S��
&���ԩIwȮL�}9�!2%baF��и��IO��/���p��5Q�n@�0���x��=@���oH9�oU��EJ�����5�wE��ˬޞ���d�U�G����^�2y<�K�.�J<�HՈ��9�*D�7)u'�ihB4B<鋳�b�l���A�E��jܲBn�TG"}\1�w��L�-�'��;�i��9Z!����� (�6ET�YZ3$<p�.�C�Z��ƍ�^T>�mj/�.'%�K�V��8��Md��_�&>f�(�YA0���g*g���LJ $W+bup�^�;���i�^R��<�~J�VIǾ,�S����衲r�h�䐬�p"-R�V�2`PQJ:�ءEAf�N�,OJ�FnKO�m*������?��&	��Kk#i �����/۔ڿ�L���jS�^��o\v�6��}��]��#V���� #�i"�?�������K�i�@�W�q�R�[L��c�(�=��p�0���I��`=ҳ4/��u(��fs=����XR/>����4y�֙�qt�1B�<�hn-Ɋc�g��N~Z%� �7�������M=i����G0���+�x�庤|~�1k���"�+�k>*͔*��0��Uv�3짞�hX;wI�s��@���N��#T�炝�?l�e�������|�8���<���D#Z�Ub��N�<����܇�vK���q�����*^��{h�W�!�I�U�5v%��ˤѩ�"�J�7.(��uE�&򄊅.�3��4�:,j�\6��r�?��8��;�ٗ��);#76�t�Gt(��5�v�_�ƽd	����[9w(�sV��Mna���)	�[���:ܭZ2}@$n@]�D��D?{9�u�g�H5��C�T�/������qC��#4Q��l��%�J�o>v����<=
���s�0�8et��Wϓm�����1WVk'sp�gi6c1�QM�0'�R9�SS�W��@�(f��甇d [�b���i�&��Z���W��>ͯ���Js&GvdV���F��Sؼ��E?h�c��I^�o��.q�%�%�gyc��{l����
��?_{�������I2��oAO�sK�JV�
pYuJ��K���a����Q�����v���	�����"3-��&��u0�" �*D`WJ���()yD��5GT
o�j�Bz���Vq�)�R ��Nn��")W�X#TC
�ly4��$��Bt
����٥��*��5^���)�w����N8�\zh^ �߮_��B���:忉��� ��3ĺ��r/�W���)�{���{�t�=Z���?<j\`��Enva=@C�xgz'��Z)�S�WmV.O���>kN3����QOQ� 2[�**B=
�pתq�u� m�`�q?ɐ����٦H(���)�S���%3#{T���mq�&�(''�}���z�z�T�ݺ���h59�ڛ����"ރ�Z��J�����n��\��񠘆|�Gv.!���lX���#9�"�����@�#%{Y���f�Z�Ka��SEB:�/���`���b��7�QO>���gb�R!�Uf,�в�$�c���x ��H���R�J�3��zu(FhwO�n�ɳ݃t�R9[�.&���-���"H�v��z-�V���"��&��7)	����Me\e䵯tc�B���
ʒ�#��T٫]�i�08���3#�gR��:���_�H>�mRB�A}�X�m'.���,��gG�Bƴ���_�2
G����]޷�L���z�~�j�P�j���N��R�<�N/�﫵�N�0�3�˝zu�m�'���)�`;��&f�̜U�e�&�����)$��#��擌���̅�3 �u�:�B=��Đ��]^�H�w�,E𧌅�b�L�B�X!ӗ1�P�h����6���2%�2����}(e��QlU�lz�,