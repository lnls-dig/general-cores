XlxV64EB    2074     a20�-3�K��l��ܐݕT\��ؑ��Ƙ�;�o<i�`A�L�ȝ^��ܾC���g�WsC� ��*�b�t��4~�Q�8Yu"b���v�y H>����!(��]�R�ރ���J�+�%r�+��!B60�w%�:\�6�ʇ��$�݂vI!�bsALH�I�֠)�D��+�[�Ņ4�*�ռ����� �O���p�'�W���3*rJ^�Jrb�����l���0�m�E���l�&`E��%b�����_����T3��b�Wy���zU�2���_�V��n������v��4{#��ǵ�!>�J[d�~�΃C�!�m��
vڛ��ΰ�x��9%��r5Y.����-��U�F�nN ��-�p|��+欖{J����񘗪��`�5&&�n�¨L_����퉺h������/�;�(4��ߚF���G��l��iD�)�MzV-ǭ"��e���p����� /�PbdmU0h�TB�֌S��b�r%�>ҟ8<}];�n�&��2[�F;��z	&o�>����L�V���荅�r(���$b�&}��IX�-f�mBm"k˃M@
QM�+�ˬC�J~4�Q@+祥�!e�.!e�Y8������)/]k2)�]Gʞ�n��l=�z���sԑ�<3�[��C�Ū�ЗWq>R1��d����NK;��?���CX�A�b���WW��)��pg�
��K�Ҙr���~(���=k:��ur�\���(2���Z ���(�=7�I3?��U��(��
^J���;E�J�5�5kk���� 飆1NV�G�U��3a��Yn�uD�	[��n��}�N�Ȕ�_� ���2�W��a�AфL��C�=�����ى��V1�!��A��yq��ԇְ/��_�]R��ƀ<��J��wSM�5`�	��?����o��ósiL�K�Ý��Q�r�E�.Vz}�3�w
w�D�����o�ᜀu�s����N�>o`�>��N2m�0���p���o6��,��vե��Z����zd\��&��J������7����1�t�lt��k����+����)#b����^VT��I�!٣X&�,����DaA˧��$�p/�mj���Ц!�\{��k=�a:Ǹ�Z����Tl�K���<�^�� }��?*���.�X`5��F{���^���P��P���bˉgt���}�Z;�d˘��2)7�j
��z�F���X��%�]#��oO*دg� w��#��~�ah����+�ӳ��o�E�a�"؆��/�D]W�?j^�~A����?��DoȪ��~�}�@gx]��l����r��)C��H��d�$�g��<��i`��𓴀9T���4�Ӗ�r
����J2F�q��0�P�)zH�+!-I�7�}���q+B���pZ���C=����(ג�����7�IaP��~#�! y��f����� �Ad�N2u��ɭ���m@��v�$����.��Z�oi�2�mHΉ!�x$��q��_yyx�w�M9R������e��S��;�� ���*�9�D��u�kc��]�1��|�vy8 ��Ę�Mm�qcv)�5~�;@�g*�K~+�1l�U��Nao���1������9G(��f�K\���B34 ��!��tki`��jZ�F����å�q�k��T���.[{�ȁ�5��7��F�����d(q�E�W`nk2B����d�Ҙ}j���w�#s��,���0��dw0Xx����\�<+��D���tcږ^�W�����(��`&>m��F�Q_y�.�O
ۘz�$��羜;b��4����)����;,dj�����ߣ���Vzũ72�qXBy��rE�9h�L��k��#����9�:Z�R�Bno?��z<��)���?��!Za��೯��9^�Gθh;�	ʡ����E(������*�5�Ej?*+`�9F����@ӓa���0|G->��<I�z�{�C @\�%��ǬP�^�Z zJ���f�z�j"?֮�|����X��2E��.����̗��c��7"� ����qa�s��@k�J6���Uv�~H�vn  �����焀Ld���؇}X�����F8cT���3�s�6�,Z�Cd��~Gbn���w�'��fK��}����!YvH�'gꟓqo^�iR3R󽏀�+�	���|��}t�L��[�S�s���~g����7��Αǣ�x5��H �JHaYP�Y$=	�QX^�75���-y�o��z�����ΰ�G�}��HL3|f��894O\˭I��g-������Ȕ=ʆGgp�ʁ�^�u{*zwOTM'x�J�W�:2�D5߮�'��Z ��^ʵX/�3�`w��ل*Kir��|���+��S�X�h@��U)���l�E>S+)n�h�W�"�-���6��+��n�Ǿd�܄��@l��|���f�p�:Ob�Nup��Ȣ�¦ao�%ZS�g��ō���/}s8��a��ˍ)��i�
��?�EH8��ߣ�pA�-O���vъ��N��