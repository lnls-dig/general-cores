XlxV64EB    4155     fd0eۖ�=e��	�Dp�<��,j�e ����3�N�����k��E�m�r@5!A]�e�zMÆ��wo{��HB�b
���ͭ����j�>��EI�6cd��r�v],��ťȁ0@~�ƍ�J÷�ٷ�S(���d�Aɐr6N��	�c�~2h��u�
�u��n��H����|�)O�ptʟ��ș]���%w��c��)W�Y�ebL]�c��(9�<2�)(��<L�>N��]�)���{+�FS|���z���b�oS���=�l:Z�^�b���8��S�a��%Z�k
��^�.JH�<8n�n���J
�Eטn���]c��=����b~Ar�W���g�_g���F���2\�6��k�$��Y��bq)�^�X��_>���3�U�ol�is��DS�iE�=O������8z�Cu��\t�nPrԌdI����}��Pl�Lx�Tl!-:׻M������/<$�����'P���x]����+�@�@�B�>�aib?g��q�%6�E%�|�x�:V��(;!�Lˋr�㢳:U�>�E�ޝ����������}JN��d�|����m�r/*�F�E�Ǐ.5�&�3:�;��,n��/4dZ|��5ɡV<���x��ԗ��I��w�$����2���}/�5��hg�BЩ�d��w��t�� !�������"�*�)��K`c�k�5:�i���݆�
{���#WT�"��<�GP.-P�{��sD_9�(ɦ��^�?B��6L������F2��+ùsV4iu9�����=B
}�x�U�qv���jD}�h�x=�����Ұ��.�6��*Ljj�u�=A�K��l�!����e�%į���>~��n �2���'ݓne6���*<�H\��Ȕu����q�A���Q%94�ټ��Q�'�{bh�f�	��K�~�~#D/�����Po�*�$rށ���4��T�K
��;I1�4�8κ����Vy�}6�,Fo����H�7��H�K8�Mu��}��,���t��۶Vx�Q���f'���о���;z[�1��e2��Rp �coƀt�P����a>3��_�s-�}�z8a;�d��%�閚5.H�N�lt��*�fr1�s��m]Z�G̦:��]��L�]���F�(^Z�-�gk?��ą<����}{���ʏ��H��(��ҝ}�L�E	�_E��0����4�h�-I�*�{��U�7�ye��^��:�%j��zS-�q�d�������5�my<�L����A���|�������eB8����wN~K�4c5[A1�2E�����<�Ƭ��(�k�[�蕸�������|oӓ<�>����'=��7��`�0I4�A�W2�G��QX�J�Dz��8�k��/"T�i�*B���d��x�f3�/�_�/R��,]IN�h>�d�H��_xܫ}�+�ȉt�,�j�>���
N2J2 �3`�/���g�l'Y�E狭�Y~p�ߴ�V��FТ�����
�����];T
G�|Tʦ�W���4���O�đj�''Hp��I�Çq`o�-�%�L=)6�x�:�+�Է,(����''�B�"�	�˕SBi��v	�LW��Q�����*�h�'�[ݦ]�q�_��SN{W�x�-Hn��#W.�b�Ֆo=�H��+ʾ���t���Z��}�7��­���H:㊫?��DEɳ�a
�]:A���~Pp¾�sh2<D���,��տ�U�UU�Gx*/4|��Z�u}�k2 Z0����)�&����?�?
���7,���e2mcJl��K;�0c�Yq���kxN�S�9=�cX�<{��C;U�S\�6@?{j�ޫ2��v\"���)O������V4�ܡG�w�}�y .B��Ͷ3��K����#�5
�a�'X�!�M�)mp��S|�xV��1\�Gm��cId��?�K���9 u���Z&Ytk3���G�X�=�6������{���x��ݽs��]��F�yBT��J}��_���d�;%�����՜��w~HN�e��<lB��Q/��u�ր�	�	A���0��V��w�-_;J����=� ~H,CE$��Ŗ�*c�Ȏ(K��2�T� �$NӪDS����D_�죮d3ט\���X�j����ޜ��v �)}��h�?6])�RW2>,])^�ۊp��V�\T�:$R��J=C���t!Tn�ߚ�|��a�թӿ{^td(��� �ݖ��q������(����7�M(Zy�o�\'I2�ap4���B�H���)ܷ��^=���=�����l-î��J،t�OP�Q���Ĵ��۷���T�-�}��w��^%��L��4�>1c��y���7
�}�p�8��}��Ҭ,Mx#@	�����k�+P{Xb����<D�������s�����2D��=� _Y�:�e��v9�x��=L�e�_�s�TЫ�pm��q�X�g�u�������6�[�٩��A����Q�y�ˎ�I�(l�{}��~�TRVʅFc����T�~����C�&���!�ɡ�(��O����K ��:�i�!���u�)��(BK[9��ВD��>0`T�ٰ�0W�̣0���_���2��i-sR�;�������p�q�%h���:��n��Oejhʘ��M">Ż���+�<%&�^���5S/k�MԾ�^�
+߂9<Ƞ����[̏�l�9����xEt9'�*�҇��9�I�k�ILJ�Ԩ�K�*��֞'4W-R�ovE��ǨíjE\A�w����əN�	;R��3��40!�M�0;� �S��/�]���F�V�R����J�N����$�~��eX���	�j*��,*8�\[��7=I��Ӝ�,6��Zp$��M���p(p:C~�� _�Q�%T��r�6=���$c���ԄSZk�XI $ٕ`s��\�;D6���u��s���&�X�0ɣ���#5I�4��as�f\��\|C�qg3LS��2����Fj�vdJ2��¯��1�ϕ$J%i5����NH)t	�P����2�l��y�p�}>/� x���-=�%7o<E���!Ҫ%M�\�c@=�Y����P�L�b�����:�/T=��~9 �blpv��e�X�z
�=�}���Bn%���ؼ>���zk
���y��6oq�.�s�1�C?�;8[��tj.�W1j�	�7�����Q2�9驝�'Ye���]_C�yk��a�U-�(b�:�w�!vnC�R�%\�Q�<�;5��(s��C�Pr/s7��a�����DgG�vV�9~�Y�)7���x~�]�
��N�����������1�8���wX�3f�D��`�nG�f��ԚM���9E���P��=�����Y�(~�7��^_��ue�9����CHJN����t9+>!�����E���*���RG�]!���ڳ�&Yk���@���^���yb�P�kY|o/�W�z���g{�C�@��<!NZ�.���rp7ß|^�"`~��Yi�B��J��)iZ�/�hw�tiE��7�T��#I4l�g�]ЪخH�2}X\a��S�������(�"3a;!G�I������7��=��J��R��D;����W=+�,�3��g��/���$�K.�[��~V0�qCGF�ʩأm���<��#+H���֚E��W	��HT *c�:|X�q��Xɩ,2�_�&J�J��;�����e��_E2�y��{M�H��%?�ӝ����/-B-�R�Gu�H����_��Wq �ị����!��q@2w�������DY(��r�~}[�o(��*��f%��f�BU�}dɧ���8�m/^�T�B3u���U ���l��*_ HG���Fj��:�sރ|F�ժ�:��A(�	�z,;�d5Hl J���!g�H�%���c��H�
��Ѐ#3�.�K�����j�D�H'�>�� 4ܶ��X7�$�#G��i�P