XlxV64EB    7892    1800���Z�<N��ͦ(�l-�p4������\gvY��������ֿd�*%�knT��f�a~¿�|}1���{�H5"s���\�L�r|��1.e�р�L	&"�����\�	�|,���Q0ۿ�7���tМg�&Z\|J��,~
e�M��4eJ����a�U҄�ă��"3�G�O��x}���D����M�۫mCY��3bS�h4��8�vr�'�׵��M�ˣlU0xWㅚ��Hf��Q�����@ !�d۲���~a@�[�-��O��</#���2��.A|�^��{*Uk�%9�|�F�δb���I��҈.�Z���Ò{B�@�(�p�}�M�m�E���x���G�ʍ��yn8���P�����*�AGM��X����W��ޗLޭ'ȵ(@�&X����H�������r	Ϫ+}���"ڋ��v��TL����$�8�R�Hx]�wһZ�0ӫ3l��D�������)׳�`�H�)��� i�?2�/_@G��k�$5��C��^'j��sn����)B.�r������<]2�и��Y˶ׅ?�d"?�\���mB
K�·�����	�K�+��_�c�y-�'����0��Wm�N�~��ߌ$\F�< �5&z*�!%ZB�z���ǢZ����.o�����s7���������� �a��U���E뼚�7�Hg-��
����:C6���OZ�'��x7V���
�D�����\f�?]��,��Y�m �:����`6E�����}zF`���_C�ܖ̛D`�6=��+Sǅ5�L�����?��%���Ш�a���t�h$k�Њ\Mȍ��믏�Ô��`W
�����J!���M^m}�� tP7�'��E�� f�k�Wy�	3��OfEf�]l��\� ���F�N�����B�E�rţ�0�[M�0�|݈�C ^�Yf	�c����	6nL���g��q>�w�C�Y1�Y���<�V�?K�_?��. J�/mE��08�V�UϷ�G2`�o�t��ϳ`��Dw�7�O�^j��7,شo�if�Z�Փ�s˰��?r�noNy��r������+�p�#���G��d�*�m���VTu�����_��$�%�"���@���9���S6� ����5��A=���x�L��Đ3�=Q�2Hj�h�����]�4��k>�lZP<���W��qo�&�+�?/8?D�J���{�j��-�"�(��^�B�Uo�}��TbiăE3�3��x�Z�1r6�<�|g!��qʬ>�˞R�R� ��a[�{kP��,��2�)�����N.�.*V��;�͎��hh��蕥�"��)	���0�W���� ���s���u�	Z�SK�W�R��+t�x�����s.�;:��(8�81:�����\�N��$	Z�GQ@�\�X�=��/�����J��-u��@0Ao9����yU�=PbND,-3�<?vJ��ۗ迹��}U *�kx��9��7\ݕw�<�H/̌Դv��,~�����SL���'�qo�%[]�r�sR9:�K�4L2e�c�@�jC��3r�.�����b���	~-�}���Q �St�4�T~5�!�ˠ��bt/1��R�X�A��sA�E��(��JB5D�j�AD�DV�L�ʵ,H૸�|��X9�=Yݚ��$��6��EC�TU�i��F�j����}*XֿU?i~��2��ݼ%#�p��I-Ҝ�4Bbaag7�4i��.ff �X]\#�e~��^�?�W��i�V�>����ã��tA稬��ǒ�n�ZE��bK��G�8�a2 h=�I'���v����!0> 2��C�	��/��n��mڵ$�W�O���HzPX6�q���^P�([u%ǃ�h�g�ħi�#xB7$��_�P��x�H^CJ��E��J?�J������-ܼ�4tÃ�k�C���>�<NTa�NP�{����;���ë��i�zI��߼���+�G��b��#�1>��CC�� ��|W�x��40�z����ya�������q���G�3~<��t�|�ū�2Y*yr�q��~�t�	��P�|b����0�%��+��ɣ��t���s�+	-�L�uP��&8��#(��fbh���nѢ*xS�i��O���f>#!�5|q%���8C3�2�+|�10��_0�u%�n�oHg5RK����������L���?f
���yB
O6ŉs��:����&�hRD�����d Lۓb�����ZIN�Q,9�m#��Z*�/�����/�l�M�Z�0�h� �����:�k�^���]�+��3L�4�!�65�+�ԃ�u�6��־���u�n���7�1eo~n�'_X�?�Y��	�c5��s���u��:*6b^���#��@G� Ҫ���aB[��&X�f#u)
��o��5����`ucK��`��EH�D��X0��]��P/j}Gj"߼h!����|b�!ɾnDqW]��'�M��	�e��`�������d��g�/�p����<�$B�L���m�5'�D���G�5?�Fp�ȃ����F�
��y��F*k�9�?��:�"svP7�Ю���� 36��±�76�2Q��Դ��3ce�<��n�P[�M[kS U2�-s��Y����q�(c~����m��pxI�A��\*Ea+Ւ EbH��[c����U�В#�1���N@���2K�?*���R�h%����D��ܚ������҄'�de���a v�Ø�/�m�Ͼ0`�9b���̕И�r���|$��5���`ܚN���A��*�6��K0쳋r(���V�N3c��5�`'��+h1p�u�gL�!���hʶg�A۹�2G¦	�X�fM�h��F	���޶���Im(���b�'�����az,_C��!�Z���A�0]fON�1-���,���{�u�r�F�RU�t�(��x�>9�w���u��ĥL��9LxL��,�̦��<�q��z�6��'b�Cjݰ~�Ai%����u���Ňl֧N�:�4�d�O~�Tt��)!!)v�J�a�������k��i��S,�yRדcg2>Q>�,T�S���]���x�����촽�p�|�p��X�krl�^��[LT��
ПU%�otl��%��� G�k�\$�ϷC��v�����&0=�~��ӡ�r��!��=$�K�u��~��x��-��ҵ��d��K`�A�;f��+��ۅgl\&7e�4���:�#Y��;�F��]J��%"�EF�5V���Wc[n�b.�p/*���v^it�H���u9��]D`��<p(o��7����[)� Lܟ�>bZ|��yN6Yp;*jJWd�$4�\K��Ր+6�2���t/GQT��j��=�hۈKW����b�B�& ���M��	��'��۱�Ȗ�-W�T�(�o���T����P�f�"&�+6�eL�B�Y�����ل��lYJ�I'�"{��2[�	UkF�N���r��z�������qZ!_�󌶦�����#��'��c��2��(���
��<'��P�tNϮ�ɲ��\5a�1���Y��7�G��.�YiQ[����S(۰9�V��uj����TQ��S����~dĖ@�� �<�51���T��)�g\�ae8���q-�-�&y���Wc�	�>[�F��<'���C�s"�3�#�5�������Z���@�j5S��z�;�4���y⏟���7e�MG�T�k;_���!|�}�܄CU!Zr�aTOC7�`S샰�1g�vrn�]���r�,?궧o}1v\����mK�Y4��J���rX"���>�Imr'\����tvt�k`�a����C9�Zb�O��m��ǣŦ��q���H'2�|��t�.���e�((�)/�&�M�_wǘ���AuY+�]*�&$!����@�ln1'��N�->�L�t�>�`$iD6��x�Z���x���dY�d-c���	�����ꊌ��\�z��v�/#�ܪ�q�J�	}Up��%eM�3t���	\ ��<�A����7
Ap�a�������EY�7
�K�𨃰�_D���;HRY���М�=P���G�J�_���"���6ʘ�����إ;SSH��o�!ڢ��.�=@�ac׬��RA�"\�_�$b�IU�Y�{�\�X�a֕Ŭ_u8|L�\K�P�m�X
̿��������(�� ab�2p�GCn|�9,����v:�g�� ՙ	ɢ�c�Wܚf�7���턉� ��`���|Y�_Q��Q���Y#^p�?�����K���SO�m�!�(��7ٿ��nf췕�	&Zj�?4�7�,[%�ڷS�6Qd��Q���F�Tj|�]�^�FI�a~�a�Y�Ӡ�����k̀�1�`�M9dz�hԼ� ��P@���F�I�(lkg���4�,$$]�0rp�P���е�� ��Q5Τ5�L��/Xx�.���Q�gP��V�r�P�1�w����q����n��#0�7=Ecw�E1Ë������S�1!�@�z'��{RvhL�Н�5�E���~kr�e��<ê���+��5��g�]�1eNE`Y0�un�9r�ù�.�"}���S�Qg�W�k��R������?ʈ&7}���F��-|���v�;�d9ƫ�|t9Ee�9���k��t/��kH���o�|��D�#VP
k�[�����=���V�.��y���t�۞JBm�K@�Ҟ�cW0�w|��w�N�8@9�⮱�)�����A������^/,���d��Y�#8>�Ew�I��3 �ќ�5*�h��(J%J�l�K/�6w
�(��|S�i�V���7�8>����&���]/�T&�9+����\��Q�*�xG*�3;�H0�2�uWp~�*���T�P�t���������C�}"�����qM�i�|#ڬs|��vW������
���I/b�uAn�>�_���^������O��t�P�����O���`o�r��_u��$.(�J�?7� z{�ⴑoY��U_���ILSf���ƺ�M���{ޔ@{��*w1WFU�c����^2� ʐ�W/rC�M� T�%��pv��'\Zn&��+	"��Y�+Z�Nȩ+�B�>�?�<�M��mb�m�.�\�ʣ��8W,�'���B��F)�G�~H�������P�[	~�?��{dߺ1{`���Z�|���PA�R(�{iށEt�����)��o���{���Ę8�1?�/Ĉe���o�[���b��Qz�(0�{��D��#����g�j��)}��V8��W�vhu8U<1�+����ed���1@k��3��=��<�?Ć���-G�BeG�s��g%�a��0�8A(�ϲ�]'I�_��L �e�
�c$���#�|q˟��)����{%~��W@Q���Ҩ���)l��7gΕ ��y[5��h(�=���{��w|����k�9�� }+:��+)�]C~�����	.��Uw}u��{cu�.��=*��,������>� ��ڇc�hkS�Qg<��m���s��sZ����XL���`A��Ce�a־�h��:B.G�T���Y!#pw��EJ�v��%<�t�f�kO��ő���i���~����@I�N�=Ѽ�ѱD�TDz��aJC����u��Q��պ�������J���u]�z)���ĳ�uDqX��`�|�ZpD�ln=d�qY*�
�='4u!E�>V_��b��<X����F1��b,v���L��#`�3p:?�,�� =���qC�QE�D�q	_=���(Ԏ���eRq�M�>�GP���N���ھKzB�
&�Q�ٛ b��TY�7��}ע�A�-����f�w�F8 w��7&,]�M!=�N�a�,Ď=�CWof���ف�.,I����
�������ȓ��Հ1�,���j���"�2�|��n����5���!�^X��#�Ȗ��4�tƒb��1?�fp�yu��%�"?���ۡ�N���5�
���H�z�X�`B[�1�(�!�4V�"�u�c�Fc8I ��rG�����~��6C�ܹ3��m���m�׫��