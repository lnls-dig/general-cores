XlxV64EB    5aed    1190���k��~�1��3�-�~RF���.�ΗH/�D���*��.ε\q$�����6��
#�A�
���f��y��c�b��35�����3���q'���!�a�%��Oи��Wj��V>�D��L�ы�X��B��`���([tPwB%�~�f4Ћ�i�g���y��8է_<g!�~�ϟǔ���3y��QOl�`�������~Ƽm�p
)��ܒE�b>m��We�4ypFמ�Eȍ��4�/PnŌ�o�<)�{g�Ah��-����G&=U�Js|g�����THi����5���u�<���.~�G�?�}:!q#�'����-|o8˽�F1��[n��XS<��!�����Z���=�a/�rtw<n��}�q �Q�>��bTʝ���+�E���f�)-�٫t�t��tp�
uCORt�^��t�юo12� ����x N�3إ��r�lt�� ���#܇��%���F��  ��-�e�|���4s-�k��y��.|�8�*�a���S�d�.��H�^�0մL��ֳ���W�(�e9���� Ol�gw�'�R�&����W+��bf��2Q �	��"�A��������m�������g��E��b���[x>�:����^z �G��%�}�}��h_�Yc�,�������ik"�<�o�a(���{U�1��^�uM͸�8jms��(
����Dé���&հBƨ����ԛ�&�����v�1�����5p��O�E(?��td<.-�Q���cJ�w�z
1N/ڿx���*��wP�Ο�L��V��&���GF�H�H�t�WO#��\�+Y�Œ��Yy{i��h�v»�#�EA��.u����O��P���6�j��M����sIlu�W��T��~$Ob|Ԫc�f2t���Τ�q��!ܼu��8$�x�A�w�**u���)z�{�,��N����Fȸ�@�c�b�PL
���N�ֿ ^ �8�}���s�
��򺩌h�ahH�>�I��Q�1U��8�_����J��4�����~簣n��l�g&��v��j��>���|b�]�o�w�%R��_�I�M��xH���!^.�Ʌҩ+�*{�t�2h�ϣ~i�OY��Q�~^���� ���3���^���}~��38��s���2)˻wgpҍS��xC5qB�����uAіd�Ӣ�WJ�w�Mz���p��FE3�29X��0��T���d��Cj3���/���`�lV�a)�K��^�@1���O��m�u��)P�<� �ٹW�İ�!N��{�"������9�2�!��Ĭ)�Hb��g�[�(&-�J�R����Lp(�%�G�WJ���)��s*��:������/���# l��>��_����Orakۍ3��wT�5j�A�b�^`XG%:VN[�2�wؖ���bGd~�?l�Y��{�U.q��u)^W���2���	-'����fXZ�8ӤB~"x9�� h��3�Z�[��Bwd��4�ޤe`)��'�j?6��`�؂X�>Q��&n5��?�?E�,$%Tb��n���"��A���a��=��UW����<u��Oꨣ��9�+����ӹ�D�ݧ|8EgW�}� ��fv�"�f^���dL
�CC�A����������\!}�fF�J�hR��w�(����H���K8�~ȍ��[c)E�8�3��=�f;����(�J�Պ�I1�P���=q��/�a�3�����uE"�X���h��ɥ��+,gz��t��O���f֘M�X�^J��kp��V�Rb~e1S1`"C����1Ɓ�.8�J%福z�]S���W������0$	Zk�}��;�mG�ս�# Zl�f�ڽ�
�Y^l��t?�)��}��gڼ�>��I�T���̯j�Ҷ�IQWpXc�GeN ��т�g���ܺQ[/�88me�y0rvi��(��
��4�*�������,.�Mm��x?�)]m���[?�`yoy�>�Z�Z���Sj����TՖ`5֜{ ��jK��E!���Rlx�XJЌp�GQƲ.R1��M�Uت	��A�xb�V蟺��W�W�eHan����[
ÿ�������gh�m��S��5�J��
�sR���ĘU6+R��X�E�^��*��e��cq�|v��F�0&NR�N��'�iA`��q*�-��.`
?�e�b�9�"MYV�M�0��a�ᱡ�j�@������ôBG-���ƭ�JV٘ �2��I�б�~�!U]��McФ����%a�j�}�`s?]�3��l-7j1Wk�RgO�v�)و��u�-p,����P�[A�L	:�o��k6�a�+��e~?8ZK�9]�d�<$�)��] Xӟ�� l@@��� �B�.�_�����.�l�e��8[����Lm�s\P*V�*�T��Sj���ٜ�n%�̄����f�n
�TY��|9~�2Rw$�,m���s��O����eF��e0 �^#a��̇T��j�,ر����L�cy���,RD��.�/6�j��j�YkR��N�- ٽ�����M�g�4�d�'pj6�b�Ѡ�&-�1s>�ƻk�i�Af�b�A�
$�N�x���w�2�K������8B���1��Fq��d�1�-�Q�� ��Á���i�҇�I��{��c�	�q��;�y-K�H@F�%�����WN�U$���R�;�hN��X�Q����:4C�qQ���:M0�������O�S�R�^�K	�t��"��tCj�Z"�5���A����\3܄�_��Z-�����(�z��N<�]�` �h:rY�H�;�>#J�\{c��'����F1XP1�%����V�۶�)�B��x6��$�l1����
�F��/_T��`&��t�����0�������7!O��b�e<�It���Ymxi�_,��<Lk�Sf60���q��:�J4,���������^w����rX��a�l�E��/�&��h�4����#�UY;�a��9r�pf6lN��k/��e���Nٸ�.�1�����8���ip����R#���ml���h���Oڿ�2��#*�?�Ŕʘ�@�X)���C�"��_�!��#|��3�C�/j�)� �P��_7��Ѥt���1f!��9Ʀ����	&�:sߕ�{�K�3��ԡ(�t'�D?���c�"��S?I�40,R���	V���]V���,��Ou] ���ܭ�Dg�f���ɹKݰC���B��A>�K�l��I�)c��g+h5��P2T�zt����j��C˕�)�.��e}�;^���R��>��q�iX��㤫d������!���Ǚ2.4�1�����5'mƐ�2~yJ�q����-��u�pa=ҋQkB׸|8���s`M�dф��R81<�s�JČ�M���1'Y��1��L���/��/�f����f�d�V=�7�(�|"ǹ�ۭrC#<��7IA���g$j������R�r*��`��{��h������d��5�����^*��a��c��G�2�d�.2.C���uV�UBȀ�A����Je;��G iv�G'@t�|�b��q#���9� FF�Fud:"<�P�&Mr,ԮP��cL��B�rDz����fm��x���Tx>�W�����kTw�x�Y�՜����Z���E�Hјe6�MF������H�[
�#z�_���?��}x��_�x�C܃ 7��1^Y;�r����IP���wr�D��郉]*X٤z���^Z8����=̙���cM(�8�#'�D"�����_U�)J���`ET[����^����~�������zd�-�{T'�zbj��o�
��R�J�p���^)�m���Q�<��$����4��D4i$��6ܸK^�<d'\�]�Ħ����1O�?c9���V��ِJO�K���Q�^λh��N�Ń��
L�4�8��,��6e}d8�5f-�����` ��Ea*�O�^>�Y'�����)��(�鯭�����m$�¹n����a����RL������睫?VX�L�aɏ,Z~�$^��$�8�
�~���rL��=�J�vj�|�h�)�s��dP=3ZK���ɶ:��QH�hlF!Jc�tn�^j�h���_	�/W*6�6Q< �#/�������޲\}Tk��ZB�D+V��l��^|�BMy@H@f����>J)�l�,��DSlq^����(���2�4+����?np���5��H�]so��;E�k�F�NV�������>�	�G
+�@�<�&g�T� ���SV`��z��b�Z����|[rё�)�Xg���MB��m��fa����H3���{k��>M�a3<��KTZ\�Y@�!��߇��ۻ�#���aǋ�*;I��޴h�[��W_��tE��s.>�+m%Q/��;2�պV��<�SZ���[e�_x�_�TC�Ss�6��ήIs̨