XlxV64EB    55fc    11f0O1*��f_�-��nc����F6zm@TT�A���ۊ��{BƲ�߷��d4Α�T��k_���o�#C�P4E��B��*eS��.m�5I��@�	M��&R�V��fŽ虔��{M(5>���X������L�M�hQ��!0���9�֧�-�V+��# m:#v�i"��E�:5��>�ZR��6_�9N8�x��jU�A��� �@By��wA��\�%�����W�WԴy��w�m[�C�ѸL�Kŵ����Z�j�"C�G%�e��w>wס����.��3L��DR����p��O�E]K�^�⹄�;wB�_.n���%n�8�*cg�̗���w`-D��>��	zX(�������A��U�3�$J7z�坄c�q��EZJ�/�ǃ�зe@�'.����S�����Voe���`��!h�Y}�b4,��=\����$�C�6��$o��'H^Q���.��{I0��guYuZ�G���$�C�<�DS�+d�^7��#sKM����PZ6�eW�j��i�i�5B��p"��ǹ�J'$�]þ�O�������N`& �GHc��w�T�[��.M8��a���|���U�)ί�b�D����p�)I��s�?�Qx��<fJ��֣U����J�bR>���BQ"��v�?�`�K�P�6���iT��������S��w,������G���t�G����b�r��֒����*�P��QAl����>(X��� ������t��C����_+���<P�8�NR�`UڎqE矿e>e w�lg�N�  ȡf�_��*#���!<�a�Gpp)�ѻQ|�M4��sybZ�S(#�GeQ�5{@m����U��%Y���u�6<�eͽ蹾��SOR&X8�>t��	m�?�I���$\��2�K޻�q����k�/�(lHf��� ڂ%2� ^$���*c^wH��q>�g�q3yǈp_�f�?_CT�F�>?���O���aTџ'�{.)5���׹��i�L�>����>���؟�!���8@��J�H��xLL*%TZ�aō���4����YS �m��ĐN��+�W���U��RC�0�gV�o�O��٨��{>d�>"�G����,WO�ב(֥�Q܇��fu�� �/����
�ûݍ�H��W;2�_~sps|ۊ��h~Պ���Q���2����"�'+^�!!��T(�ju�\� �ʿ�<��P}�1�-��4�x�k���pҧ;`z�S�s-	�3Q�Jnt���顁D�����l~^f��,�#,v�Â�9���+�m�R?�!)���>�V��UN�;_oi�}4���Y6�uE��+�0A���[l�͙��sQo���/��EIt�L��n�h�k���+�~S�P����|��"*ڐ�o�:��q������pr2�Np��D7.�]�B�����TгgKZ���(�O���T�Ke�zƫ�a1xt���cw�f�4��+�=�!]v 3B�"o�*dqe�:�7��So��Q҄�.��e�nC_3�'�w02��x�&��t5��w ~����_RY[��{�^���3�:�-���y�v߲���-�f��+ g�I:�%�.2x�Xr*���H]�4G��M���L�&���*HCә�.��!��o�.[l��.��]�$�����e\�����z e����<�g��Y�ʕ�j���{m�|���D�4���!�ˎqٶ�	�m�����7�X��rQ�����<��@l���O���wz`~7��T�ב�?KJ��;B�ϖ�t)(O}��V�4���"k|�	xҐz�޹7Й�ԅ�$.-�Q���~��{z��ս�趰��G(�A��ғ�1����Q���,T��v�4i~�f/§vm�*5�h�[%��Z�yъ�~d�P��3#�� T��b[�bB���i1J�'%��W@}��.ʐ�n1_�	:�� ��mϫ�96/��O�ABr�4:�n< }�|�/�N}�	8�k$Wn���ۮ/�6m(%�w��X{����ש���[���v�E{�y��'��|�9��E<"ȼ��!f�?$�\��W�`��䵆K� ͇X-HW����f�>�VI�Usn�����d
�����^#�t`��4'&��#]���7�mi-��>/M����5!�ޤ�p�!��)�RLdM�ygO*�����m9�N�ڇfk����r��lE-S�P~ASg��u�:����kw��4C	N��zޚT�fFW�y��9���Ĝ�\�
�L�6��6<0�¼�F���*
�x��`ߐ�t�1�>|JE ��|5�۰x�VF�̑f՟�v�8E���G�|^6U�c��s��զ�|��4�kY�9r��2	+ȸ�����j���r�dZ�4��~�"�_��%z"R4q�	�>i=����d��<:C�E������YC����
�O|W�z�z�����0�D��i��m^S�Ky,R��F"�R�e(���"��_��w����e��;h@��	�UF��Ǚ�L|��Zi]5l1O¢>/���&D߃x��k�֑�׮��;Z���8�Tk�_�9�{���h�I{��E!
��̖�Q��qE��]��@L�j�Y��׀� �-�����٧�ȁv)@�׵��y9���F".y����YNT�qb�G{���c|<�b�K�u��N����Nw J���������6��=C��~I+@Yp�1-f�j��74���9�ڐ`�g�͍���0Q�
c��M���S,M��#F������.��˗���s$���ro��U�� �('����'FkOU�5e,u���'�O�z{��ε���~*�[��9*#P=��%΋9zѺK�e��Y������mh�5o���'���XR� ؙ����nr�[M{	���]M�l��З�7��T!s��O�3���	��j�l6S�|O�����!�D �}�B[,�ZK�S���u�|vN3��5�#�VhdO���}(<��+G�"t��N]�K��:���#+���c��Sj��Ǭ|��4�-�����U��̐9k;WJQjA��q��ۃo�����}�\$O�э���#r89Au��J�.�C�4~�i9[�.D��H�z��r(̺d�
����[��0�q��Ӹ%��R*��п����zד�|@Jn�Pہ�A#G~�w����Ჵs���+q����;���J-�B��ё�Ȕ��0ǈi���'��p��6�V�d�P�6�NuA�����J�q�R�g/lS�L�Q�gӂ�EY�-P�QB�c4�� 	q������l��g�sA���o�K�;E�h��MO�S���%M��O�P����1}�4�;��Z����h���t�9j��-i9�o�n��>��"BqZVE��4�B(���܇����mj+�̌i�� g5Ch�@�1po�q�-�F�)H~�2��z�n1��Ϸ*�޺�q��b�mE3Wy1Vf>^���#D
ќj1��}ld��>��Y��h��v�]�]�;���A�P��1�8Ŋ��v�����֙м���s*���^W�Ʒn',��pC<W?� �&h\h!�cǦ�hZ�[�I<�$����[ګrZO�˟�!�ov9�{��b�7� 5�Sd�adn�n�M��~zM�ߦv�%�� O�6�΂���լlL�H2f�.��v	џ����(�_��p����pF{��L�MJY�f�p���5�V���]'ć�ِ�-������JM-�������ܭM�Pt�M�f�+-����H*"^<$�X�X¼؛&,�ɵ����ȅb���XcZ����I�c/�H��%s ��ֈO4N۫-0�iņ���auY�K�VX\E����0q����1���g��,x��_ `P/b�c8�ʬ�h�E1���-Eek�rL)��pH�6��*��E Ko�`Z4�+1�!�i�h�3zL��'��a�a�Fw�e�x�!�^���E0�'�%l�U̀S�\z�[�S��Tk��n"f�</��V"ҙr��/k� ���=�H�J�|Y�����Ϫ�|��~J563"!�F�a���Qo!�z�G�3�w��[����	m���Yh��[��O���(�/R�, ���E�ޟ풩� �p��_`��וl�!:�5� ��O������D
�=T��i��>|;	P��)�z~>��\�=z#3w�'9t���?��|�a�h3�9S
����Gu$�]�_��ll���1����������W�C��R���3���Ib�l�����j��dz�T��XOo9�<��j�\� �AʈWcܐf��W�arrGA���� �YXe{��H<w�j��0w��F7�^��P��l��P��ͧ�	��z��q|3�;������#C+��'j�d��@��*�,{J���t���ό��@���E��H�]�?�~~]�sw븁i%�X	\�E�*S�5;��Tb�'�o�ea����c|a�{