XlxV64EB    4ad5    1050�x�_!O"�����H� �y��As8�F��7��ָ�ؖ�%�юz�_Oz���
�����K3�!T%Ը���DpG��%��:�=Ey*Z/�#��c醾a�Q���V���� ^� ԙM������) �R����w�N�o`W�O�f�:%wH�lQ%���I��U��$�,s�n�����`�?F�R[M�����[+FO�R���|m?>�<�<"� �.V�pv7��ν��I-�(�*x��+�x��MIH���,$wHr7�����׉�BW���1�D�rY[��s��20�/"X��������B(v���#N��Á�L�!!
o�IIp[\T/�F�V���}K���l��n4<���Ro��(�.�i�4!�5J�Fs�sdsTc^�J�ʂ�7w�I$�������� �e�R�5�k:�Z V�3fX�f�'����d���G���w�ϖ`��
�we���)01d��A��"�J��l��ge����j�q7>x��Y���B+>��q_���n�0�ާ[D�B�_��0�Q��1�(���&z���X=�^&�w&� W�#��b�C�!�RW���^���ȷH�I@�Gn�3�\��������ϥQ�15>-ç0����5>F�O��o�!����$u�'��(j\r��*����,h��פ	-��6��o��uu1l�$�o)���E�\&���͛ow�� ڀ�:�Z�q�7Bëw_'nG��/w�o�C'ɇ��#�d���.�}��i���/Nh&�>���E�G�I� ]�O�����=������Ա�]x6�S����.]I���]Npc�>�6�B�eE��Pg1ΫB���]�>��O�k���v�����P�l�T�����D� �A#���۰�b*�)�S
[ ���~ꩥ1J�e�D����xo�u��uVO���`��u��)eG�1��%���1��ڻG_�����I�Rp������^�a�X�@��5U�|�/�k�m�HJ�vJ	����U[V`�l���x|�Ûu�Vvz"��$�M�����)����-Yi��|��ؖ����JI����}���'%��:VN-��c�ǎ����P+8"�����G�-=9<p{���E�/X���^��_n���8���|��
������3ő�;������4�NC�'LA?f�=*Z�a�����9E�l�ք�^�c<���f��9�
���p�3s�W�q�wT�,��"_�b��m�"����z2��O�[E8��)�%��K�y��r���n��ڣ�8V#���w��|e�K g�ˈ}��/x�8�� �~I����>#˳�ǚ���mT��`b=�5��@~[�Hhl�*ϼ�k��Sݝ��w*.�gnB�(���������=Mr�@�y\������c�R��|��g�{/�Ԅ����}1�,5�����h�n6	�ס���rn��s#E��y�@��CȰÃ8?��K%�|H������⁲��Q���Hڤ���_̌���e�&�a���!�i�p�)�+wS���{�Dة#k-�����sc���w���]�%#9�c^��d�E�K����|�O���ۑS]�븺��E���.���,"��7��=,��`�_
z�i[zԨ�O6W��YD3�t+؟��T�pp��꜒�&T���@���ѵ����*� K&Mg������2� ��um��q��R[L�-*�cЬ&Y�j3�iP.���#!����(d��61�e���z��o��3�{Sr�����N_I����:Q���d��7�o� S!_�7�%)\,>Z��$��_���X��
�t+XY�^��\�2	�U��%H�C"��B�=���ZJ�ܑ:�:
}��u��'[L�Z��`��+�0�
*bp�=�ӤV�z�+Y.���dc��2*�njA����z���85`�2u��+���o亩CN0/�!S�V|�U\?�C$~=Q�k+�|Õ�IE!a���y�,:<�y��OcQ�9,3� ϲH��>��A	-�����^����Zv������ֱ೾��R��
�>k"�d��;�V��B�r骟��#]YԄ#ZI������Ȟ�T�������W+'d��x���s77)Zwd�͞�y&�@T_���|��Sn�	�ê`~�<��r(ӧ������sۊ���x}f�����A~�M�ӳ�U=J&~�؜J�.���,����@ɤij��S�iK� �:߅y�$�a�d�f���ƾ�S�r�
I��/� �{e��b;�E��:U�AI��U����N/6#o���4����5pd&#Ѩ�9x�(į��zl��,L�w鰵�_.��@2.OF FvZI��"&@{�WDra���z�{�Pk��|L��4PԢӥ�8ۚFr�`�\1�X�**&e���	d�vݱ���U
�4a��"�O�X�;wज�z�����\�}e����}�
{��Hw��K쯱S���t���{%u-ۖ�T�$?�c�k�/\�Rx�Fzȑ�׃�t0Mow!o\k���Q�\)�sE��	���A=Cm6sR)��ך��|�<Rc�J��Τ��0z�iDy+Z¤�5s���$��f�g��%o�5E��"�� �����c���p������S������%7])OTm�+]����;�@L�\��
�u'KcN�:o�}��I�K����]C/r$2AN�U�7~�O6K�"��'�����'�ҀőB[��w��駫���[G�o�Ϻj��UX���*�f��2�c��GQs+L��W���`[������0�a�8~o�8��d�N�-�,�ǆW0�S�2X�S�>�D2��1�S&�]o@6J?P����6s��[���{OLý�x���xg�an�3���C��n�������a}La
���ۢ�\���M���)������/�g�k��/C���>)�(�:3�	���V�/kp�O8c�v����Y�{�.���P��}�G�|�hA�?$��6�t��,~/��6JU<O�i���;�W�U���3���m�5�bK'u@L�W�?��pd�%���qh��`����9c�K����;��N�j���g4�8+<rIf�ȇ�mT���^�n��p��c����I��ʥ]���$�Z�9�"F'!���@Oœ�i1��IGR�&��.�yy�K]˨�X;Jd�����W����W��%��(����:yd���g�?�q�mc]9�"C��Z��Ev���ٴ��*Z��N����EL"��Q��oʌ'7�Yǭ�65q�
h�Ī#_;����|��ʶ�&��o�8�Xc9	w�V�N�)J�Zr|�@�/��D_�*i��d�2�U�[� ��X�G��Z離N��A�+��l@(�^�:�w��Plφu��ML��Xw�� f`�e7���R+,�	�Z�<��<��D�s����;ΙC��cUsK�6����e�x��P�0��Z�F)�$�=�^��X�Km��ϲۖA	�作�-����UDg.zӈ���,�zR-����x��_�L;%�؋2�q�j�C�>-ts\"-��O��c�M���~Uq{f?���Ci�M=}�7�u>'J�1�D�twep K�T��rT !P�h�ӹ����%Ԧ�m��"��=��0��|�-����.�y���cRUK=50�Ķ�us�
Ql_]4����Y�������Fڂgm�y�t� ~c��n�ޮ�V��$ɗy�[K�G�͌�:m��A]���>�4�ti�Ae��$�T��\&y�	����E�M��j��4tǖ�K!`x���f�H��G�q�Pֶꙴ�s�8��0�҅�8KHa�z�2�'�/L��G����v���_rxhJkd�'r���o&��Y��(��p*�4�uDj��?ҽ�)(�nǙc����~�6E#|P^ܩ�6m�1S�Mu�	��,6��;�%2jdt���$W�S0�h3��RÇc`;�OPfT]�FԢj�@����Ap��Mq�	x�A8�ݗ-�7_G��!�M���3P��<F�)&�m���@R
Ê�������l�>��Lzٙe�5(�C�N��E�$6��^��"T}���