XlxV64EB    fa00    2480"��*���D7�� �	L&�@��ػ5BiQӽ�>6k>�8ы�Ͽq���j��Y����:�(����N����ѽ-�7���G���ݽ����ĺ�Y�q��tP�_�F�M� ��fe�`<6V~B��'r��ĩ����\�hޥΡBY0��Y�JC5;�?���tDAC�>R/�puк�������D���A�IE_
���Ʒ���b�G�T<�B\�k2/CB�
����c���%���ޱ�0D���P�h�)#�#V�)�>":G:t.��(����>x�<&K�t3Ř��Ң�k����an�+�%и
�rd\�O؈8�ֱ�|��/V-����l�Eӻ� և�зZd���0w��̉��W�3=��/������8su=Hʕ���:�/wH�9*�^8�G_�|n�v.Y�=��h.�S�s7O�����ؿ�n�+g�ѣ���8@��^u\]�̋��sd�]�����z��3����i�/S��Y��B��(�:��Cf��I����J,��Q��h��PI;^솈��}&�!� �
�c��~�E3n���Ŏ��xUT�II���M{&���n-�p��m>Yў�&>�ȸ����U-}����J�sD�D^opj˳�B��]ܻqc�)nv��Ϻ��Y�����:�����q�O�����;N�ʏ)I������̀x٧�(�`���ΈZ��#�sf��a�&]b}���۱���N������?/Y��MZ]�<��U��Ymk��X�u����g$*o�y���@�a�z�>�ʖ0bG���߲��m v��s=橝���[�b\t';�e\�oe���F��xOx�4U��
cdj���_7��I{d5��
| ϊv��y,)�y{O$�����c�	!�qE�`=�E�p�J�l����k���x1]g�Ď��U�He\vK~���X���	W�̇��e��0�'�J���کi�e��JJ,%2�0/�g�γ �l#X�B�DԌ3N�h8hL^::�����J���a 8�֊8�wY��伀�8
�s�SWw�ЕevS�(��=�_��MVHY�^=�еc�yka��L�o��7sz�NJ͊s�Yt[�I����u��$\�7beӫK� :Yv!1+�?r�]��y�.Г'������� ��>��w0}��N��������H\�X�y�����u�,?���P���߰�׮`2���[����R�({�4T�������FN�N]v5�4��FO������EIȉ���5���a��D(We����(�ۢ�m-^*�%g���G�*��oL�=�`�������-��7�I�ε*VD�p���K�L�4��Wҍ]��Ѷ�=塕v���ZA�{��o�_��X$���q+Q���:k�Nq�!���b�' ��\�Ś�vAڅC�'�L?vt��>W��o�x�x��:E�v9:*�s��g�"��y�с@���1��:5�z�\`������o�E&�X �ӹAz߲�V��U{�z��(5��w�{��х�1��?Ul��E�ˣ�-8�Z��f	]��\�@a�8P���ρp��O�Й)l8���|S��p�����2�7j�3��F�<��Y��%3H������iX�譐��}E�)G	m���;��JkW���� 9��_�����Ax<�c�˕�$��� �%I���q*8g��'ˑ:�ᘘ8�yJeDǓl�R�z#O߾
��b@��6���*PeX�nC�k�E=����������d�[F����sL��=�$Nɶ�����s�.�?������g���~+n�16��h���F$���;ٴ"MIH�h[uc�C<[�*@q&)r��sD��ڀ���P�P����ȝ]/[�������B�5�k3����a]b"0F�W�(�j�x�=���&�K�{(��>��AW*�:qΛa#㉗@����j��
#=�W,�8DEB]�N�D���
�5z���E�b�(�v�/4V�,��\�y嶚���XɆ��b�Q���|3��Ii{7�|��7>��(j���
����Oy1f�4�)��Y������){g��"���٢-Q/�u�&�c���P�Mx)��U2o��E�U��>:�8�.�[q��Ba�3$����s���鲢�C�F&	<f�a!4&@�Sڧ���{{�����[4�0���r7��F�
�+f!�`�")�m⃽5�LfG��U�4A�l}(�7{�ʗ�P�|�\Tpg�r����5`���ʋ��zs��:5����ι;g֜����I8A�퀖��6.gR�,��\�%n���2�ɧ"�ݰHq���������㚣�j%�6K�'��U��c��,��~<�X'>���I�(%�R|[?������x��\�Tf�����Qg��=������9���(Ҳ��`*�kU'�:���!�^Xy�.��|u����N�ږ�U��j��s#����ȫ����X�,i��#��콣x�۔X�#�c�P�<�9�s�gX�=�%�Rr�h}s-�p>{����6U3�J�~* �/�1�>G:ګ$�`�����Pt�!"Bq,���<��E���PaN�AՉ�3�u��ty~�ܙ�^�Hijv�l��
���B/��#�#\�#�<��+hQ��A?�ݹ��$�g���҅=]��(sM�Ի��*ES.�720�*�eV�靅q�7��HDz�>]���]�hHw2XA�*&�ʚ�z*+��Zp�
ً��h�d���j�6M
,�J�2F�������<*GMi)�E/���=�L�����v���L�*Rj��Eۯ��I2�K��+8؈�hʂ�T	���Ëm�U�ߖ�����"��ƾէP�Ñ�!>�*�nh�����'�|� ���w1s�`g�3/]����*�m����A�c�{�b��
���ڠ;�����?SsiD�̘����7�8�������$�V}�rP��)���8l���ռ<�FVw���>���9+>�gz��o&��Ũ��d�G��؄\�$�5ٮQ��a��q�yW�nx��fm�dt,X��
K�@�#.��1d�޶ r�GDI�'x)zz�]�6���e��b�P@�T,�2L���߻x���"�ܤ��Q���8E���XEU�;�y����ǔ��z������x�M�
�ܩn��ퟓ{$�M����^��G]T=�S���/CIþg�!Բ����}�s���� �_�g�"�$�hJ�9�7��"���1�Kj����Ļ;"��_��$����*�3t~�F�e�ףD��_9_��l�r��>��0Q�X��ʬ$�S��O.:m��4d.�7p�X��ɾ׳J����K��Y��9��P{;q=ա�3�flV$�O)ea�I�>�niTVH�j�>��L2�M�����"~cEj���D�~�ab����QMoYH�s~��KD_	׊�R��wb&%����_����Q0�R�����j�x�­�-+�Ju|�')|`�,nT�40�����EA�O������ɕ��쯁�R=�̞A�H;f!�����͞�o��2ۈm�����?gU
�/B��ʞA���Qv�0�#\��n��x�]��:׻#����]���6��e�	������8�
��2 |��)tNz��p���lŴ�Q1TUޖ�Wq��8��m�6�jX�]�Z��@���w�b�����4���b+S5�����M)e)cANG��'c�96�0W$U�pH&����$"�7�f��/v}�����+;2z��X���X��<F)��-�|4�^�g�S�?3�.E����vb�S��@��%0'�<�6*\���p����D��#�aK�QE���ʉF�%�z�C�3A�]i4����E����x����"��[7�%S�K�Q<�5�� ��
�9>�yu�8ӢF��ڲ��_��2��:�)���xn�OÊ�� [��������D0_#q�s:� V�ZF������뚨�`��4S�wXl���d��z$y�+�m�M{��d�X�%�<BA�cmE���~�J&(�w@0=Y!mv�(t�$S��:�v���h���F��ނ,��p��g��7붠Un�PpAPL�c^5��(V��2,K���y�_�{j�b	X�������Ϫ.����8Hz��?�F5A�I��Z���E3亶��E!iV"�l ��k��^�(�r'��EZ�{��qݸ��P��=�@�[K%d]�Xg1��ZTlu���ϕI1��@R�A��	�_�^Y��X|�CT�`{Фyw����C��0��Cο.�7 �|�A~4�`�lhh�y��G/
x��r��j������#:�T�_"��Н�k�&Š��|�[D-�ٟ'���D����z^\c�p�~�1cYY��W��.n}���QWZ�U�q���t�n�:tZLXD��¥G"�%�gL�S��#�,u(1fQ
n����qs�����y��~��S,\����3���XBc��@E��o���� ����5��8Ⱥa���@����>��������$���%�ۥz��ܦ1��,���Lm��u$�l�A�*�"�;V�e�I��i��N8*)*T�m@��X>N�[��vu�)�͂	��vh���G��N��Q_�O6OI`��2~��푖�V���;j�rf�`�!E'��`Է�2��.7�ë�rE��D���G�L�>P�o7��%�i��i'��ǺQI�+qoʺ�N<x������e�5_m�쀖X,�:Eȓ�0�I�0?��z�oM��f@�:ێy4�&Ջ/PI�,@��j73p��}��J�>��aKK�<�Q+f0:��xPJx����5��;wY��<ď�ٌ��L�v�����Q��~O�����q��C���=�s,�@p��� L��[G#�}`��`Ƃ��s~���7��AÀ߇y��0_BTY��\j��_ ����=��i_��mwV�}��a!�v������
V���0�Qϫ�D2��ڋ�(�XdQ*��C[l�>�;�U���c���;洔! iɖJ���]1߫��d[�z}O�1�hϊ=o~PXȟ�73#���儠	��1Y�v��������bW�p1��o�r՘�wP�4W_�,ِ������I��ƃ��xp?�J��vЗ�2�X�8.5�!2�gC6:�q^<��U- Ҝ�ztr1���K��?(�Lէ\>_�^�=(�œ��X3�.Ƥ#��z8�+�"��e���� kW2+��e�/N�I�"�SIy�詘�e�D�`'��ܪI���P�u�Z\�t��#�U�c�M5gn'L6�e�!�:��a�κ�N��\�[fՏa�6A�;y��P��$9^���4#oT�G�2߽֩�}��3&�Y��o��Q�����i��if�X�#K��R5� }^�=���Xu{�Խ�!��7Z�
[~&�� K*��
�sĄL؟z�,�cqU��E��[۽F���\d�-v�Y��N�.K�A�:5�x�=�g]�� �`tU~�H��^5~|�C��ub��\Z*x�a�7�JvH]�\����%WB�j�zQPdQ�xs���3�n�yL�<�⊠G��G��Z�/"&/�~;�'��iO�������V���{:�S��>����DWa��]Z,^]�h��.10'P�e,����j������me3�-�M>�Ƚ����>�8o�nqK0b+X�
v�*��J\����+����f���5��-n��P���Vn�%4(��pb�����vS��Җ
6�;<?��/�R~�f��9#�ə�PO-�[�%����0O��������{Q�+��� ��~j�&i>�H��b�/$�ho� �=��8��"03�	 �����U=�������f�� �4�`�V5�@��:d�&( ��$��
�(�!�R���fOzn�,�W��U�G�wwO�hTm���F�]33�0ðyl��k��o�����Y�����*�Ƿr�&F��">�.��.F�rN����1T�+7[ȴ�S�
��)Y�]|0j";FR[9�S4=Xhr��.�P}�v}
������c�ɖv~��`ý���k���8hYU֓x@C��${k-Ch�}������x�̋�t�ֈb�K���>a�M5Y�P�F��W=g�$!���Nm���� ��˲	ۻ��zm��!�u�[�n�W U׉��A���1aR�sX�N�C�gCrɅ��Ge�~3����E��5Nf+2qJD��[s7`��1��/wϻ�:k�6F����!F��>�G|`4򭔐��v]h=<����\]�	�:(#WN�_�ܯcɸ �������7��������� �kV�C�X*ܟ�[�>c�#��?˞5�h��cQ{�l:}�m��QpT������� �)��SJ�@�5��m�r!���L)���J�=��,j�&}q�M�<!#�@s|�v��+,��f^�S�Go�X��kt����<�B������=USW|�`���RlNB����Kl	��o�j��/R%�sN,ػ!���׷8�M�9�r��o�;��!3E6�%�o���8���[��b�Q�De�}L�2G�Gtf3d���j�
�G�"A�bF�b�p��2���ށzgN2�
��P~h.�������dG7�l6��S%���g����:�h:��L�P.�FϨE��.�"�'��Y�ψ!1TD�J2	�2�ݐ�n��s�^�^*"Ll�U欧��mu����g$��Z�IуQ���j�_������p:C�?��B�d�hR�����A����lr���,lv8���N�7}����]��10B���rF̡m����x�R�[�.�S	�ٶ�l�s���F�؝xBFg�ʩr�ܳ-�= |����e$]6�^#��/�]06��>gT+b�Bq�
|J8v
K��}��@Xβҧ2�x�J�M�A��θ���O	��t�V�㗼�W��������霪��H�71jW�C/��~�=]>���'��3LFy��1#��1K�0��h)V���߇�g7%!���� ���PSU�9K1���q`2�W[�E 󛴗F�͈P��=�;�F�)�|0���hgXUZf���������É����j�v��wvds[�����P�Vtp�^���a"8��7�+P�v~��L=��б���������}f"��*�z�'�T�E�  ^Z=Ǹ��]'���G�19���B溁9�*年���v+�u�����(��:@��F��sz�p�G�����0n�z���R`��0�$ezr���C�\���[�*{��̐���f� �*���Ӽ{�K�gn �Ƴg���օ6uSpVf���5�2W&&P;dWH/�!b4O`�� �O��E(�E���ؿ>�yҐQ�PWjS�����/P��d���7ǔ���o!��� �07s�p�?˳�w]�2�|1GK�nQ�������z7���/!^���^�X�0����lJ��Q��V���7��2�X�W�xU�4mss7ݫ�K]�iP��v�"�)M_��9�e*b^��� �e�E���f"}psQ�N5�%�,�#NH6h���s��d��5�m�l#�&m�P����K�4,����-T1�m�XGLF��}�BF|�wB��X{`nf�')s�ǐ�]�[#|��c�;;ʬ4����k%n�H1�'F��k������ܝy����"�״�P���c�RpX��T]��Fa��r+t����Ǔ�$�O�㯅�*��QdE)�4+�zL����S`����'�Q�����.�u� ��k�(\Ĩ��V�l=ZdL�,CH��JB� ~V!�8���J���^�nq��Q��K�@a Lf�VP��ָO��m[~��b���F}��>�t�n��\�t�T�5j�!��O�2w������Tj��J\�J6���| 3���x,����h�]�A���b�N���5ܒ蝗�5�vRa�?l~�u� �bykP||b��o�1
��k�F�'�<��a��*�δ{d�և0����W��A >�_>қ�5���H���t�L�/hpMUv�Z9a�J�V�ECOݘ���W]�r���}4۸B4�/5]u�ː�Daܺ_��z���ЋF�~��S�1
1�'�批f�кƽ̪� p:�����Fǽ�8O�v��=�]/�,M�:�|�����R��.��	�X��״��z�>���
��:��؏���9P��˃�j�b�p�S*xA��B�ik�P��Ts���v�M¿�9�HS���N���:Bw3\�Ȗխ���U�q�L�t�������o��d8�\pu��TA�`Ō�ab-�3�����x!�-2�����^�Op����6*�I��"�f��.L^��EH�c���g���IM���fc�,��!+C�ҋ���׮����j�;���w��$m�]��$�~��&��5��0�	�h�&mh��10F��m
X�P�	��{��`KtO�4��l�K�N1l��46��D��=�%��Y��&�a/�1���'/c9.y~YcP�К����¡7yt����'�����AaW���3�( ן��;oy���{��h��W¤�w��Ǒ�,wJ�F��S/ª�s�y�	'��)��S�]�d���Gú��f��=�+>r΁H���T�q�N�Ok}�͠�x��j��09�H�2�*�����@�^���Ԝ}�&��EC��F���ˣ?��B�Q��l��56�I'�G��'��"7�`�e�3M�h:ٸ`u�,Q�e��oyW�쁛�B��*7K����Wi/M�42>T�
�p nbH}
yu2�./�x�"p����T-&+U��v�m��^;q�^K\��El���)�y�i���P"L�$�5I�=?��O��)���:��I
�@�\� -M,B��:�O�DYX6���:�1D���V�j;k}�+n��`�J-����2j)���يF��t�zI��ùF�7{0y��-�������P��Z��W���4�1F���O鍚ˑ1pI�d7�6��E6@SX��7��������h�����x��-�o����d�/%�A��N��-&�^���oP�F����;�N3���D�|�+�j?����Z�u�;�^ff��;����T!N�̦�b��5j��yr �+!��ϑ�J?h�:��c+t�y�2XlxV64EB    a5fb    14d0fT�E�6r��,WK�˩�y������?���w�?�[7n
�[D�5z���L�v��v���n-�� un���q"�'�O��>��
?S�9/��H�a7(��Fx:�U�"�}�PY�dz��$85579�Q9uR�=f�9�5h���Վ",���p�R�}J7	�U�,�h�&�p7�A�G��hIW���Z�Hg��+쏕�<�t� %�)+�t�H�
��. �TXefD8*�?����^� �S��jЈ�`ū���|�ط�_�:���]����0�+��WI:�4ߛ+�P�Ɖ�";�9a?��/�b]:�3.�ʴg�����������*�#8lR*�g�A��g�!Ṗ�/�C�!?�Z�"���9NZnLJV��wI-�C�����=�vW"��P�m|^��1��=�9�E�Y�-�N_�;i�	�\��&�&�B�ܙ��������kA)\O|y����S9K.�X�1^��Tm�#��d�`n�0��h7�����l�Y\�5O�
;"�=�AD�gJ:C�Ep�ը[3�,<��� �O0��]I�ޟF�<�����h;����֣�E�3�~l4]���z �3]��7::��*N��lZ��w]����	��'�������S븴����[uεZ���ֺ��+j΁:Ы_�b�/g����ī|��!1�{^ 1d������|uZ�^��F���H����S�ZY�	|�x>GPRߢ�s�8�K:FA�EΨ!?��=X����T�@�Ra��`")�8�5ݮ�b$�<����.�Ok,��xzS�BjYF�����(�T2k�R�4و�D�8�!c�/�N[s��Thߥ5_ :M5��i:>�\|�k���1�&�a�I�7�!cGHP�f	@S#�-B�[`{v��ld��.��/�� @�NcW��멉6lY�6sdn6��c�'OwF`�t��K�u�U��M�-	M~wD|g�)�\:���m)>w�T��y��&g>�VSR ڋ@u#�L�l��b�����=���`U��_�'{KA���t�)s��]V4ãS�:��X[C���|������εv����7.rӢ��{���85&�D//�C��"�Mѩ�a�y�@S�]�hs*�z�S�U�PH#�5�!�(H�)�m���s$���Oٴ4��忦��kM4�,A
�������LU|i���8]p����B��MD6���od\��G*��X���-(�[pˬ(�S�z7�!�bۼ�8'ً�[J��.Gnc邻Hdkp�����m&�Ꞻ8��֨�'aĤ�+��Q$�~Ðu/�´��z�Mk���Ռ�+���(k��,�-��/j��"u9�kx�ú�]�
z��ӂ�'61/���,��k���]!��X���6�c����@[���# Ύ_��@��;{��]�}2Y�u��0͕�=��jZ��Lv��	��[gF����xz'�es�Ne3��ҵ��|;�	O�}�~����X���Ť�'�=U۶I�X��݅.��I�w������(�$(>'��8
5ś`���7�+�T���Fk�;�*4��Wy"�����m3�G�<�z���AM}S':;9Qc���_��~j��U&~�k�����&����T�)��}�vo��9u�5�St��{�r���-��F(��j�_��A��Xk��W�,U������
V45g���h��3 +3�L'��(������,��=����t���s�Y>4m
�
���e�/�"�q�ɦTC�
��<�F�#e��~U���~�U�@�Z�5���iM�Y��=�]�����.����������AL�K�>|�e�S����g�35j�6�Mh]��ѴS5�&��L��ӊW�x�Kp�dj	��4�L�I}0���L|r�>}�㽎���G�3�ʔ�����,���]��l��| �56J����ˉ&}�o8�>C-U1�m�2�[4I��&Ki���R�%�奴����,�r�0����\Ãl�ZؕV!VP>ee�^i~}j�X�
���D� �Ռ+%~�� �m�B�}�a�����xO@�)�~���뻃�P�_0�62Z_��L�>*��Ϊɛ�X����>��
����JU����@ݨ0�i��n��H��9Pz�Ov����1Z�~�B�L���!ֳ^E�]�B���R>����]؈�2��`�
�E\����dݖ�hzu.yRG�Y��5����%�9;��W5�C�a��e�H`<ʂ\�±m.���j:�ܽ =�����ŝ��bI?�7����~��%N������'�v��*�ÔYnT�����E�'�7e'̈6�s�DB/y2�yl�ݱ�{D�	�<���7�"e�<�Fq}U�m�.6'`���ypʨ���Y(�+R2�}b�g�{�~T�k�D*�&1t��jwb'M�����X"'4�wdN%G�F��l�n
KR5a�IY3�&��hXxI"����Υah��١�wN�����TU�{ރGpF�!A�m��>��o��ٟfbW^Л����#�:ޘX$��*��@;д���\����@�h�v.���$UJ�P�1��+�Mc~�&m�W��O���~�B���N� N�U8�����]c�%&_������4�J[u�9��X-,�}&#����6OI����>*���fc�B��M��F�o��P��F���/#@^���(`��Wh�?;�����L�6h7h{\�u�_V	F�9��a<EGFyL:��s�Hs�A��!�O��Ub����x���h{�#�.ҹ���E�,�y?2�\�Ȭ�i4��RW�`��]nMZX�P�c�4�1�W�G�jae1��"s�C2.� N�"��N�x�Z���Ϯ���ؿ�j}�{ez $3ƿM}"e^h�3Ii�7TP�E��Q�<.d$ߏ���>��� 5FR��Ƽ�����~[f�!z���4��g�H�W�89I���
��YhC����'��I?��$���?�|ٷ���L��R>��ȶsKZ��J�^t�ؙ�q��S�>�V�~�z��H��pA$^�5��3�X@r�`@Br��K���=K��:W���tq>?%&��^��O-�j�O�0�2�`Gb���d#��*B��:����op��^x]������q4��H���$�y�J�f���;}��EB�6���`��q�s�o��5�oyT4�!�Ir���f9��1�����m�,u��Oґ(D�$��g�AՀ>��hXb���Ӂ[��;МGN<�~�ɯՄ��{��Q��耟i�U#,5��4Q4�<�f��q�o0���cg�I�T�#�An	���o;�Ƙ���H�I�\�%�9[D�L w��acf�㹎��� �Ve�]��l�Ka9n�o2ú�G�ü��C�zT7i�5�Q�n%�{_�$��uZ����~��9h��& 6����� �2"����l����eܮ<*lރM�l�9��	5ZU�8�&'HV�'�����K�<��r�c���+�u R)��>:�xr�`k��b#�i�R����	���[p◴�9���!J��`�ko^�б�����j���&�c��/z��H�F2+琡�Rn�ղWo��-������V �
/y�����f�Ym���36�aU�J{DI��P��ba@K�r�@����qWI+SxYݒx��k�m}�- g��]�k��wK%\׷�	�M�d:����Q�jw�{�ͺv��+7O8�!x�0oLX`�qp�.Јt���
����D;�RiK����/n�:�j�l:?D�@��*�����E��W-�
B� -£p�Px͏��x5Rq�a��xW��0io��;2�$�:��;��6���`Q6Խ_������}���0�ݿ���*�u��	��e:�:nޏ5qV|�D�3�ࡼ�S�c����s��U�L�\��O��e��u4�%��ڇ:pcA/8��W [���=��W��6�'H�w����A����a��lc<��Ʊ^���&������"�BVI8�5T�{W�(Ex러�Q�uEIȻ���$u��4�O��5H/Q��k�1^��mSII6�8��Z��rKqֹ��_��Cj���"�.�n��������%kQ>}�4lsv���E������/��BZ\M�2�H�Yϫc��0�R�"xf�1ɡ�x�7.�5��3�pyU�y��U���WB��F�B��j�vį�b�!�T�%��=�K�����a�����9@	'�i~�*<N�%􄫸�h�!�1t��l�ZEq�qo��E��������4�<�]a���.̰{��V�����#��5n�q��;7th1on@;��O�#6�#TU�����S&<K�:�"�CΊƈ�-����/��Ԑ?�'KN�]���ɍ��b$�� e_[S�{zװ?�����i�5���e��� �?ă'*�Hו��Z�L�׻�ۣ��u�p��뜬�)�\�}�����"���E_KP�6\�x�IP���ֳ�rS��Ԣ�EI�|��F��|����(��A�Iv4\�Un��r^���}�.xn�ʗ��0���˿�%�s@���CM��=-
XC�p����S�A]Nć߲��i�Ý�W�U��nE��Q�
���\ӄ/�;$Qht��ɨJ����~Fkh@
�(��XMڟ}m���=�K��0r�jxv�e�$I�E@Po�����O�F&�ʗv-6uO&Ne����Q��C?^� ��{�O.��TG���I�}��3k2Pu}�rR΁�	��|����<�]��9����H�!\T��f4Dkp��υ�o#\���-h(�z�s=^�Px� 	���Lb�0Vϛxb����u����6��ta$��2�+��C��V��������C�U�*�>_�}�/���s�;V�����$����N>��)Zd�m$�)��Ι�%.�I���MK�W�`=ώ�KN߭2P�OqO�S����N`��,U4���V�-��DK�*���Qz�����yX��a�u#,#�?�Q*�������6�\�l�u��M�_�,����[���{�I�?r�X�h�k��Ec�"��h�/����d#�4d ��1����`x���8���$�&x2�l�%�;_��~��앉������m��o�XT�4ٱ9]-��l�/I���C�"HO������@��ަB5� �6��A�'mr�G{��T�gzk�1O�/�O