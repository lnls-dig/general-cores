XlxV64EB    1a2b     8b0 z݌�N�� k�c�|�է̋����/ê�`���+0&[�w��ɖ�D��u�}J���6��+#�0,Q�']k��[��yB׽��H��5�k�0�3��i�R�\No�Ie�h��P䝪��D4DE�>���SH�]�]5n5`�E��!�p�jf�XϟX����}{�#����p|Sj�a)��P��������.ܦ=:�H���kj�5���W�0�*�"�9�>m���sgJ��z��}�N��M�Њ�cOf�v��/�_� �]�@��ȡΚ����9��a��*[�%�l[��;l��8e��eG:=�o&x�9�������W���B�y�x�ªyeh��eo��{dtN��>��]'>W�j������
��H
�rExWXo�!l9��l�Kt��ȥ/���z�%����K�K͒��q"��5d:���f�9��,4�t�u��l��^��j�r)�Ո8��1,�5��j�ڟ����7!�$8�4�]���b�R�v,�g�j:0,O����衿d�y�v�B�Wqety"��ђ:���#V�!��O�	I,��d�|k�~�kp��BƯ���e�J�-�a���i&���r6];g�XgL�̑��gd�u{m�vuQ�FK�x�,� �_�9��ާdsA��S���ǬJ��\v3�RkSֵ�c�J�f�����~ Z���7�h꣡��V�|ҕ5���X�8],��4�B�2�nU�#��w,_�k��J���������EJ(z�:
Xr��`e�Q6��� �>i�9=��$l�A��nJ��3��Sޢ?� GSAzG��/T}{��)MN0��M���!|}�����M\}�`nc�W*
kƞe���If��>����si����΁�c�`&�z,T��:�t H��Aǡ��w�#�����]h��N��0%�I
��j����W��(�Z��>5��&8�=���:�ZC�z3ߏES&���X-��JcЀ���V�
r��ٛ�9+2du��l��Br��p&֌��g�4�D������/fp��_/S6�}aIU�7�	��,U\���������cOm}�ȹ�P?�@ƤyD^�lz1�2GuQ���<Z	'��e�㠷��N�S ���{*,�ok��:Tr]:�>���9,=��)�Z80}S����I��²j�۷؅ޔL�UZ��	���V�v�;>���V&s��
[��p�~T�MSZ_����,u�Vi;����x�NZ���=��c:����>�Eƌ[�p������m�ϸ�e��)���q�W)��0�������/�x���&D���3DP@GOF��%�����4�#���L�m7j��ݻ4D]���=���2Dvف������<�u[N��3奺2h��E�ą���F �i��t&VޔqO>G��t礸�r��⠏p&�;��L_k���=�[e<��Z�[��?aBA�E|��ɳF�͖�tB���Mi"�:�8�=�.tn���/��֭WC��1\	q�m�c�!��YƓ���v��ѥ����9%���9��&�hN$��\u�V ]�B6����W3zM�-5n�AO���^̒�ϲ��l�ԛPb�N ���r��n�"�-�S�j�J���Ht�u��{>�Qq�_�v��{�
H�mG �S�ܤt�%ۤ@E�^��d�1\9ۂ��.�2q)Z��"mSVF��b���0R؟�v/�����Oo#q��l&��{"U���3KX���?o"�R�����4����`*hK/=�����|�M)�u��"��`Xc���|ѭ�`�br��#�Y�Ww������0r�<+!�A����!�
3H�wjЯ�R�����������}�C/���� k}\.&d�AF���1��4�ko 7}���e0.%��-������RO˶T��v��^n��.j7��dB6.g�N����]�z%�=N;;W�g��	�m�Ŋn? �hzAT��o  ���	&�K�'kx&B���2��Q�0	Ϥ�0|�c,0vn��������-[6cZ�,�?"�,���T�㜫<�e�������{�����T��J�1���$I�w�F!��5SN���{y}�5���2���)�8V�`���"�G��	�Ӌq���(��P>^hL�L�Rtv��GY��O�V�1��U�/N ��@j7
�H��&�=�w~�֥�G ���d�