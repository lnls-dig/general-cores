XlxV64EB    1410     7c0[�"���hN�td0,i!����_܁h,+�c��M%$='�tk%u�?N}�����r"�]j2B#�������({b�2�9���EӒS�d��ݓ�^l{'��C��n`2���H���qf(�p�k:�I
p�5s�}����E[��w]��r�R��΄��r5�!��Q�l�a���wx���`z�\}�=Q�q���^�u��a�ZU�wJ�2�|s+L��ߤ��s�Y��<Pe��}N���oO6��G��}o�i��/�>$�}�j��n=��y��*\���a���|nzd|5��xz�r���u)�]�����N�����'d�^�S��_�Ѓ��Gz�o44C��'S���q[��2Cϱ�P���`�2�xÉ{pރ�x1H��i��k��[։� �tP�Q��8@��gyC�Fv�pఢUmB���ë́��҂DK�E2�^i��xʹ�_$rJ�0����d��;�Ѩ �1�����o��:{AB�Dt�P3j ���(j�^��0Р.�-�O����F �&�������>vr6�G�<��v??msܣO�!MC��F��z7�B���!%������U�l���`LwN��f�kȕ��\��&n���M�:��C>�>G�W�8��sTC���G�|6��W8�O9l
��F{�R<���/��Bg2{=�V���\y>�6��.�Z%���|�}���RO�9��nȲ��-e\�K�K���v�{���jXO�I�-�"!��fT8A��I�Gz>���fd���Q��� OĀT�8��*�\
�0��ͺ>�&iQ3O��w��ﯡ���/\T�w���b��ɬX}1�oq���OF��vq.������j!6���Uf)�u��V�T-�!����7y�+1�t�<B~��	�N�����f������Iu�Q�u��f�E|���A3��)ˍ��P�"o)�WZ��4E8((j�PV���������G>���ɬ0�S9�U&7���;'?U�L�aV��`�IT%�i5��#�nu*����~�mW�Y�skE@GVw�-Y�݃��]�Y"�y���:�ӣe���ܞ�D���o��!"���%�І��(�Xm�P:;�t�sj��AO�3a��)�d��dH�(�a1�Ϊ[c38E|�J@ߦ?���m�悒�����L�m�o��ә�D)�B��:'�)kr	��ke]��A�!���m�o(��C��-��du�Veޫ��lz�~
(���r_d����de'��6����<�#��S�P�B��$9����D�.�h&�M�� P���$��������o�tgo'�yLO!�N8^�-'Yl�R�H��R����0�����:�W����[���̖uн��oD��r�J��?������ڞCw��L�OL1�B���A���M�܂p�-ǜc��Ȇ.lK��]h�1�or�����m�-]OG�l�$�_���P~ЗC,fa�x� ܱO�[YO�w�s��Tta$�=y;� I1G
�{��U�UӅ�ZI&hQ���.��	�$B5��/;ψ�COB6| fܒol�%3���_�>C�����ѦZ��9�0�E6�J�D�m_�U��ࢇ�u#��K��Đi,�]`%.���ERmQ8b,���}���6���쭼�܋
��8T!�J��୴!�?W�j�LE)���䵔�ۺ��e\Ƚ�2Y�������=����1��ț�:9T $��Bd:>ص�^?t���M����y3"�EOA�1��%���u �ߪd���잡�_	�^-����)�N�P?�j�if{G̩E�:`���m1��i7d��
�s����M�o��'}&J-�:�AL;���bU�rP��5���H%L�z5���O��Bh�rڇx���QBN�o[�&���@[Q��$��X�`��n���ˋ❔,�a��RZ